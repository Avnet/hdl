`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
N5tpJKQsbMBmnk3gnbOYpEgbQ8e5U2wFGmjnUOxYsC9tZe9qpuCGTN7BTMmPGuuaQSFSWzVQ2F/g
9EHL8WG2dw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pPWgujFwklYtXX6kdLC19fBEwvxa+l4hvV6hoET0ylSadfraoYle6mRuRag1ouBs3DiTA9csg2X/
3OwQuMQMCL6fHLWuhuID3j/8/xfOlpBqRrC3pFn5GdPdCnu1qgzN4ps++mvCJVvf0PZppKlJSpaQ
BK83L1Vdqu4Ryul7W3k=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vbtWWyNWIgvbYDUz4JCNVcAI8n/IojqjjJ6DSQPBsgWS7JVLdM6tHBD2JhwsDPjIIxdMvB606Fs0
dwTkCrydWMs1N8MYzGs+4ErKcMkW644gMytpBaUiJz3yzJHJlOiL3NapCjPJ1q1WSPArzfA/N2/h
CeRXlxUPPtm8EH1UcNPADvyUPu11lhtNGJsdz89cjNj+E+AFtprV0phM9V88LdWvMIo+DFhu6jF6
lssQJd1LqUxeZuXzfiVmg7c+xO/v9LMY1aYTj1WbEpVK2oEEFfwxwO+AQ7rADwqv3LduiyWw8Hs8
La65fjGSMF6nZ3FoRwLRnANaW71s5wupYsXhBg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KMlX981wHsPDKOrJzQ4BSXb8F/2zAqIZgRiA0dyhUS7DON4rSCEyvGQ9qsdNAqjrNfJIkCRhkdkG
Ktx1zmgx95Exs2o9N7qTMNvVuhQl4DkjpGZbHsXpLGcLicVZMHyFCNX5RRKe26cePpV3+VI1ICwn
Ok1cA/IWTbcUJ0/6fUIjd4K8s98F6MoCkf2OFDifBzg5CFOpR7CrU8nRdBG8eMOSrIhj+DFdZfYV
cqJWxTp2SIakQerljVJM4HMyechvkJZdwOzuI7B1xSo+Evq4q58EtyVH1btZt0YydprjKMB2YBS1
1QdF6GU1bFD8Yu4ilesPOHGvUKscu+Vhxu000g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ViM/4BCtDAxGu4oFXi0myys7AvGFRqQxMxPdWM8YXNConLPjHNxJTKP9yH5wazC02aKAaEUwA9kg
7ltfP+Ee3M5N40XjzAoJLhv1kx1kBO2eRlAzq9J/S4vahmInF01wo3d8++24BC5fpHdgfU3SIs3R
ky1jUQOkim8faV395jA=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WxDi/+P4p4PItgr5nEP8MI4kjQpUpYpPHJBzwl0/RXSgMyagFvd1KcmoUVn6lZ6QLcavy4MZR2bX
zhDUyLqeBzO/UkssweOxBq9MxdzfQrSS+Rb1qV6LsqWrdQDyuMk3Qzcoez1FuhOHYRlMZfZt/5Kj
qn6st03RY58g9+Em81R+uCG43EngWi8WWEgd3fJ4ezx6qmaO+kXuWSQpjHCuE+rnnGPHNYUfBM5X
9Lz5mLMHBEGImjkYT0GUmtZn7MXinu692eD/WiH+CnDeD5hTMrOQhAHbbubJjdg7mwHjeyK9YpuB
aTSKpsnKfQ6nKX0sT6umtahK9FGVCjJSm89D1g==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3QoWuftDZmvyfRhFgboz42YjSObxF+eeMBqD2lTWQV1J035/rtjKm5Gk6R8paoGS8Q8QnhTLgJAl
rl/zRIUI+ZRdPKwAH8gjRYgYoEWYU6Pu2SsL4rYIUo6ilhRMaE+TWttfpeXtehiVL5h7yKLS3BsC
3NtrL6uQPTw6rab16yZBEUtkv2tBjMJWSH4Bv1Zgi/eKdNa4/XkELMtgU/vt04zSHNN58sBj9qMU
aFz0JODSzNG4tUteWT34rvB+FfSRgVhXmM7Rwi2nubCKVOoeq9N07ypQx3nwnUaDX+zaUU/qNzku
IVeah1Z5+3Hp76tA6LbCM9whDIA1iuaXIppTdA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qlWbfVLllNsKIdtoZUi6ldNUWRYS4uLr6oCEXay6EFkdB2HpwSyO7NmyczHv7J9qK4g6lTDoRhcM
5XZMNdyK8bvwYmvtgRWAihTLtnsZ6p8b4fv6Wri2BwwXS7fhc7/e3f8D2lHp6tpsgjabJNryNgK5
xlTj+bgv07Oj2gx/WbeEUWqWMSc8zth09QsdvDjdl1GEIx2mu3xyXXfMXxf3rLmLmFbjvpp+xk8R
AkOB+TnCxpo1j8OPzyrmkcw41GhucRjoLT3Zif2LAavKmUZ2DaepcHc3xgEiiPlhxDetJkiMPZdp
rYvSDomBbMATOTrzfWard2/Hhlsx+ek9u8eZsQ==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Bp2FKHl/ru2qBGFe1nS/b39yES/r9xQhrmcJVr2BBeBbtU9G3EXymrGKxnQSsE+bcybBgbCcl45d
0JakwNs6vBuS8mvCA96jNDuspDX7LBYV7wMMwDGR2YuGVA7AtlCEN+9PrE3+75++mOGOjDjO6u32
Pj5Unl3bMvYDUMj4R2CNV+bLkFsWB2cXueIP1jUqsIy6kgFMLoMX4vAFFu+J9GW2hJ/CWNDMLvdg
kRKODhfeZk2ERhtiJdOLWxapUGQP6N0HKIOuMuUPfzGi6gwBpLVyYpZYCfkKiHTxZM+lQEGqpBJn
LavYPRXndPyxGxNLbWr6y9fgNNQpetFeEaj3Uw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 868896)
`protect data_block
x6y2881loG0ZfSvZtu/jFRjAxEDvIjKHRXkdk+bzLctVhyZPB28b7N2H032CNcb4lpk4vjc8i5AA
LXaxe1JetlP17KlukVBqnrC/vgspuhsGauIp+C65j9XlCYlZuIkJDrsMsTem6eBgnsANN8wmvI7r
fGgUYT8oA0oQpaAfqXfD17BS7+AlEtCsb8Z5+/Jyfdhd0N/laiOYRRKnH9zEC7UAjZywxz0NFbp2
5Dman1j/z6E1CUR2fpSyI/FjnJXTycw/3d7EEb1e7Mg2BQ703uWXqCyhBNqFWihcA27Dl7TPQB9Z
E9IQebYQrjxW9whyaOkROnew8bHXri6CUui0LTKSIWdEcZa3nnDyVNM1CYVzSutUajQgPJ2wZSiM
nnTPo+4BcScXHcAUbjCcnkAEhYfDcyWldlcAPznvdJqwxQgQ3yIMaFYifRV6S4mCczUh6Zd4Hi4F
vh/AqfeJ4iI/a5aTY1ZOctKT8zI+GOQP91UiRtdVT7gsHXeCM0eZfT7rFCo4DnDS4k0Csgz+rj06
nnZ+WnJuWFe34Av9VMSpOV5eB4CGwtNDhoIRCRz/h6xLSnEEl9PB6ydjWxnGmMnz0YUt2Ytnuwrk
zPdp3J2iQZZhle0MIucima+PVfzIJmah98UjKcr3wBVDtja86ar8yz0y8e7UJU/vhtyHl6FRraJS
iy/aASFAg2zVCsqB8Ub5PAWDIH8B/vN0GtQSFTMcGg+74dbXqIWXc8BQYrO6M+zeNHRq/vyJC+Kn
yxMZH70DCvlfTs0+Z/lK8IqB6Gnq6hKP3gWzMOO3wejWGPL8lXffCS7PXnoGm2OEAQmHPIm7SQaw
+S+sv6RK3L60Wu70njp2exMns1g8GKx8KNdKv8E/qnPGoFst4Y+njBrGcT7CeczGEQyyAA3z1SjD
VMSpM8jm6KIsL7cQvejA7ojjSglmMnuiunbBiRC6yEQF34zBOsQ4PygudNWxRn6dJmOs28+8Fk44
OU4NrNqJoIZyRorJq1gmknznJZKE0EuzglI0RGi7JeTR0lOe9nxXDkgmr8i91XxygA1iV6W6u7S0
g3pTDM6fSt6TEv9VTcGQvgJ+k1soHC5MN2NNUDoQAo7r9H7uebxVnsqnuYt4bT2AtQw7zUHh2e7m
kv+GQ5TB8aefKa+QBJbWnxooae+VY3RXPy2As+9PgLKIXAmyFsm7QILAE6oVlLZS8s+aHgn3kelZ
7cSOnePmF13TNM6TjMpxYKatCvn+cEYNQdKeLptHAcnnnxp0QJCiRsS737rVtaRudIf1NvXXD55e
r2Yxm7RXBQ3KzFiE2C2DTpLy+gGScgOprAxcb2mYO6JFJOrYffofszuOJw4YuWfkOBdNpchzlBNq
qIkLdeS4DwMeoLDvyt3/NhQlR39ivESZf7vQBn7xPDF4QVmk0XBg5/APM8GzUvNRZMNFynWDqUX/
I7m6R8ufujUSIt0hnWDdayR9Tg5GdcteFfGM7F4x97badrmkYi5cwpCAcUFMCPdHPx2+eTRJTDMb
HJCxhEFUauZ8GcOjwqCm+K16izoQYXwamzLXBw/MRiywE93hNN2NKG5acmTHdEeFN8seTXamWxMu
p1UBADV8yuDbPwjt8yZHJQ8+OOo/lNlFeR/qk8OylVGSm9/9vRpzpRHs0x5bLYZIJOm5uo48c2IK
FpsumP/7NFOhp5EBoTIDJCy9Sx7DzSjAhGstHlWPcugtT9+U4+hHAEsXnfAV9KLOq8Hg9ruWOb9p
sgLRN8YzUgVCckYbYEkeujQdzDuHQlAstczwvlQW+2HdH6brjDHUQLgwqfo3nLHjqjiQO5ib1PKl
pj0F0Fzz0E8sxZF62Iue64E4uVTThoBAdzhYY8O+1VST+003hR39CnsZjylVK34FGyNY4fKziisr
GZQc4ALXRgTZawvnpv2YFeW61535hiiUwblNEcgSIA/5NrfFeOaaZZz4mR49gix+yGuJgyocrhYZ
s38eD/gG7N1MAP8LUwAJb2K2iPDHBREmtaPXg4psl8noYWSWJM2ScQhQ4B8uJ3gYbCI0Pl5Cc5K7
qTBhjLVGCbyHq4gP/gEeQ73tv8XSc8fAT2KuxmaZdx4nKxxhIJDNgXSCPjV2dRvlHqQILlJxWF8l
im4OzBRB2IA4ujVUPbCBy/Q+aFtAEHTO34o8gTfsLH4MpkjxgsMOJfdQ6ezij2xcdSsnc/F+KNUj
HKubovmPWhPeSS5aWjlo8MLwlAd7lFlV9JE/hs8Q+42kpkoejjL5Lk8mjpRDeqLKry7j+Qt4uXPM
PCIQR3FFTXmZ9am+pNiqk096JzJzEj3sxbwgLIEzkgE9zjjWpDn4B+bvmd/cjC6q9Oaz3AXP3gy5
lOHHGNX0bQg+OdawE+2ubFadYBgdOl4K7wucEhN7Z+2g5SXqxRci3Kbiv9dkyQbHqLFjb2F/NVOF
sqfdocMadULu4pBVFyQr6zcXJLiN7vD9cmY3T77M666/KjPeXZTpxBz7UfgDr1wPU2TOdxDNiIXC
vbPBq5M+JcvOhvBKvhTulXQGsMnmLZSWXth7VB4vTTiPjelWUWxAkHcVI4wOLdjpmPed3xOX8Z8V
Cm5v69hU+JbdALiBJ1xEYbrkrEKBXTdobJUnzrJ4JazG2/zXxUvJXcHAp4LH0hoXE3bTIwoyNHB/
gC6rsXqhnCLHADgCpMuF73gVEay3OZ76z2E2XR36HyzLnGan1dvJuwYr/zl2SJqRsIyjrVRGBJGs
dZ/oVH55nptbSC3jLMGRKjITxintBz2Gsf2EClvrN2gyD2PadnDEoa5TZLe70NnmHY3Zx9jelxyl
KLLTyP8sC3SBMn09aoe0dvqG9Int1ODOl2iJHboJoZaUQCtJHCqOTySpoqG+k93r44C9YfQ4kGkf
IqetEFY9Be6t/fOVf8/dwEf5/KQwYZ7KvWAze209IdgedX85Wt6HI7Dm8///lPtHR/JAF6S7JWIY
wdx2VEr/LcrX+YpGCN6RrYJ6dUDkd5sKanF20PHnivgmKqIinwKNF5Tg/Kavd0OGelVXGSmWO9L/
ceq2pQ7C+lz3LDeUg2UljDiXC2dsWdU4gIfH7qRJHivbPizP7Ya8SdRMiQxDQbXzJWQkA3Bl31/m
EAGEVcuRMiPA6Tf9GOqx4uCp7L1VZpOoSWYEJCBNYlHTXitsSX3mm+Rn2wQ5r5LA2nDurTfHStr1
jbv1UL5yIRrqk2a8IYLnEkJiNUHVStSzfyn+g0jY83Etj7oEunkd5Vy0CaoY8l9iUK3vqTdsetAc
oA89aXfpnXyyaddcRk46g2E6yUNEeKyzOeScJRd8btMGW/hZJTJAlubPDpJ2fyNUAwEbF5xx4QnV
5abcq06JQKUKB9y6i6P4beZpWEV7Gi4EsN05IASedCrNIlyHLrJhfGRJoLmijmPqOxRyaWINjQoG
UGuJ3oQtXNr8RviMwH6SBWFUAEcBLLKq70JXvUzbOH6fpRh6XB88kxtFC4B2v0njWL9SX8Wa6ylI
X14dCBEGCJrg0F5GkWVxr77dOXOsBUTc2/uuSycj7sQnggIxfhvTIiVV7EG7aMETBGnc20zzfiTT
rWT+37p6UmK4FX4i7SqTPo5QgC3bcZedrn1OdODfDpjFFtSR+g7Qvoy5OKexA2uhXi83hCGRQEwa
aKpWRi2E1L+tKraro0xP1b0L/1RwYhOOKWbnXYoD7pa5I8SGvPu9T6mrE7vz0TYluUx0n+L1UkNS
AiRz8uvuiYac0AFLCb08fVRHoBmCT10vrtFNZSASfcglsvOBnDX/3O5yYJ+N6HQagg2EwfuxchBx
NGHlA6oexY5acAKQNQu84eXxr7SwtyJA+/gM22Ao+TVb8QtYjHLelqzhyDlh/hrp63jEERUubOb8
CS2SY0/6uqhPqPw9YV6ovMaLPqxZptSgzQUtbtt8fpDw4OojHd4iH9FgWUFsK6M1FAXe02fPmY+c
LSyu5SaiT7AMom54SO05xJOikpCqe7PDxTwT7rPczDSdjvXaB4j6VzodexLFjv5r2WeNSCmzYTYb
nqRuAQbfcsfWnfWfE5SVgBeiwJfAynTL/GpJN7jjpgwqCjf7oLA/9AJNy8GLNotVYK0zu0XnsDOw
b7FCXqDuEEc0RJrAzezaw6ZZI4y8MrfxoHAwiyGIwWZz/J7cYGx05RGavxfjSvvOE2zcJVf3Li8u
PF8IoHUgxn0hX/ve08Kt6aGQdHu13G6RWL1nxJRVdk76zlGkbBa7Q2KAuzew3Z46m5NH9sy8hOGM
/pjjYFDCWNs+y6cfAXHQV65EcqjsrRE6c+SGQR53PLDPQMhIBYXyH1nPUg9vFiMLoFYwqkzkC6nh
oxUvlkx9gAnwB7L0j3vPp/UQkAWHRRYiGmHpFlNtxDlFvQaFLZcrPsZ5EWhqesAAA63+mo0KpJyz
yiNHigz6jnlxKcLYiDttxQhxL4BYrtOfDRqFJmEgf2zLEyzxj9Nq4c3KIG8s8RXs4kSn4buxOY1X
JzUnR42ekP+DpGr/quX8vgTgg4hBGbI0YgREcEr1u0wy95Y3T0BHeyN8aDgqz40hVC7Cs3PZE/ld
C2JLeCDGv7+8GmRaHFSP43ACL0SLGWu8x9FprAjg+J/7+ULzePmyWVC5YfUQR/iNNCckL/At8Qc0
oxwTy80fyv/4EMR0r64FHDzTgKRl9f3mkdrfrFmiGiTMMlrMC29L1eBXTmOWnnAfRqdpKcQo6m9f
lV87YcE/gxTptxnXvib/0NMrhzqzhhBCUaTwd9OZw1J1GNhj8Dh1aBnU0/Qr8AuQDizDfp8nV7AF
lrLXfZaEHSRFQ+uUZTj0egqxZsr5w8H9fhcUv3xxZE9S/t/YHMlaTC4LUtYcLdmY4FGqttJZRhec
kIwMbaRxw5vpxwafwypNysqOQFUndpOBwy/W/2pXg+IuScjJYGtNGUkxw6g1pxNUTcZ0X5wRxuBp
VwooeTOhuQ0al3Q8b7vSNFPT+vBmJOyK6Uojrdl53s4GX7XxTm+CckbC6kgaFZUoZgyX7tFEtndN
/4sNKSHRRwILBQa1UYfFAMv2d9lwlmmbgYkG0PPADoAJ4ZUUsoH21eK2M2xESFSt7F/cWfysvk4v
s4Ub0PNvkhl1TuQTTpqJsh4kjrJ7mBeXMQ7huLE0oKhMvk70yPYDkmxdOJLIj9TcGTByzbrubfUA
1rMEa9u/SSj1FOk2DlWTh6sYubEkAZ2evWUlZ/h4Q7LJyAWbmd6W+vcV+/Gsow9/BNEqdjUOwdgt
/kzQzAU9ye6PDEnQNN4H5yDZRyaLfz+wqFO4xfiHuGJbuWp4f0x53G3d6vYzxhiFx/EsuntHNI2p
xQX/bhJsh3rl/vp/6fyE78Dt6/X1UexvhcHSPaNLCSUYh8oMLsZB4XpkmSRLc4yEvrLgGinQLbEu
FCf0goVLy5HFPydkL242oH3/LySdCnf8EPbC267Oibozv0jiAITalIwBho8TNrEsHYEznXoWfJGo
oebO2SP9L81wJ4xnmDc5cvtyastFM13Rp6kRYhUqjSxWsV+bjfOcGuxi+JtL+9GnLfyoyArgk3W7
FtulzYTG6ac181cI8oStJbu6g2q4DGWeTZlFR3gKtWp3HtawszhQNom8nPeNtXC+6HfUxmmLSuPC
gC+f6OSojE6+mVyJdchuJpKCRPMDb6MNhNmRPwVipT+uK4l/uALKMnvBBU1BLg8He8weiaE82NbB
plhjN5XA+k9XWUBhsu1zZTLHUhTLNuB91mVPsy+w0KhBgHphudoXd/OXOblsFXb+mREzsNpQcb6o
8GFTqlakGJJAAIXLn29KUpORy4WPuL6sTF01Cn548x8+cI8gEGiLHqy67iBh7djqN8WLl1E3Mt2h
RDejmDXnWGw667ZmyCH0upoTVIkTaB7I0mj6zptyLhEGhx6KDh3NLMW2Z3gNIfGjNt7tUCO42aOd
MYSyJO6I8/+B0RpQwt8yxVlRWVZoHzuQTA0u7Qne6IVa6bvNpRg2n2JtN1VPwC0X2sCWvj9RZwtf
UF7teaBKuecSwU9qfjCSp5Sw/QNwX60SnD+/+SybSZwkEQd5sidIgrjzJZLUFT80vM+nWaUm3GTF
C4MbbLv9nrANXcJX4lhPeWo8oUq2eDHMTe1FIT8HJ67nVeilJOY07p1KnpkajP3ldE8QDm+9GFJb
+Vv6IOaYCcSYzMDKQgPvGIg4HgQ6G6AdqCV7YNz9Tk8eqtqZQnORP9e/CSLo6enx0TCJ9H+LaaVj
Oi9gImsvqAxfR3z885iH4xdfZDYLkGZ0bUwpTtpCfwowsStjwGsN9oIw6+y4mdDz5zb2KInUdIML
FA4lA+XgAC4poCIFMmZVnecHfPpcM3FLeneZK51RiqMz5LRg7Jv1CENTJoIOMzdyCEjtj7W0oiXU
4bxnPZMFTq49kTAcRw1psVwpwuWHHgiDFkUzeSr3y6ShLlQlIRmKCtM/1vw46CTFEa/21IqFflNw
LOtKNr9+ySO9BGjDAHWKd3zO8QbkQJUFTFJ5AOL6Dew9DdRYOSNMumW4GZ98WPYFFI38wRMGj4Ta
9H3/sOwsClv7tv5ckO/Gac3RSiWJNBfKJxWqNqZew2TQvFuESEqcxArsFcQ0wpaAmUOTaywCS/Zi
4JhU2U9+t2mw/nbHBfI9WEAzs68h7qu1vxH1xxcU3ldwi8+SBaCoRMFLL0Fbe7jbbcUG8JfXrfdM
s8E98gEjFNRtSt6c5wZ5x5wAQZn9uvvyIVyYlhHsBx21pwMe+3kgqQ8O7u4n8399T4E1ABXvG6Es
Lb5AH99Aowd3ZHq5M8yb6DIV6qMviBm+KpdWJZ6mPAiDFb9E7/pFIrwGIO3bYfKqkitGjm7rtX0y
gNQIW1MPLmXSZ42alGJwTcLFuzvtC4exGS/ANy3r+M660j76brv0Iuv474Sg408b2NQKcj3FjdTN
KtiGSbPG0LYmGfDSkdMo9AjPEI2FXRQhShodUwjqOalGtq/4IXj6gYOt7IdvUTJRg6SZYDZqv+56
zkXeMzRpo+468LVbMGjBpxyurVEn8eWF57inQIc3DL5F2dplKax4dTLoCkFoySa8TbtW3naomgqt
vMrwknhuVMtZQhne1rXh9VRGvhtKvv6jMl1pL83ujvDokEaU1H/sWi4/JoJnqBiLzpgkCWaLWbvh
HbTdzzAk22nX0XHUqQFALum+lVucDVJfjbi/rlgqibCAVuVMAkLNJuUMaZRF4LPV1mSh8xmOIEpR
8EMwIDaCzLBWUGfxUbMLBp//YoJ1f+1geAirLaCdO5r/r5sD7OZw/RAXf/yPJyiUP44s1Ym2buDc
lGuWiCp3lebOpfwxWaozxJJl4+pMoEz9EToSO7Mny6Yc3ArxfYaxfXfIQ1xuJByGHOIa3pBG7B5X
HaM3uTpOYtvx4tlLtrK48c70rorFaOiSk8VD/WOem9fJPIGcwqvIeNqCNIUEzaLYbvczXdam3h20
AjX4tMtN+LzeR5QDPLjS4bC6OVsbZv75o3r8NQseCe8obXMue+HBPrphHzUo1UmxVEhPM30jvKXk
Ui9RNCbNTX8bnz6BZIJU1K1mbTrctq/Dy97BxbiR0JH4oDOG4K0dx944KBSN3oRVFgq7IE27XwjY
shSXmLFGiZCDlyQwp0OQ9ZUIu5ZJ6L3vPBwF94BBfbVQkCdFwHO7ijVSXLOZQdzkeYUkpkZIBe9r
KWbvSnWW9OF3T60eL8FyZCgvCdUdKt3hsaGmxgPnGoVPtTxE2BSioYReyMNbUJg3IzXcPBYodLTu
1XJ8uynhZxivh6EnNoWWAhyZwx680/Ylq77I8TzcoSSVcZ/vzBU5JwP16FVm9dYyDTwIXi922wPS
sP9R3CqD+GcwzUFRdBunz9xosWpU1T98E08bijqEIy5lDX51RC6XuKpyi5ppHP/CluZi4Bk/Jxik
bGPCf15iSDOkn+ki536Fxla8uIEw5qj2O3AtyU/CzbwP3xuoEZqUPn7lcr8zOegYTw4/nQQqQFqz
cIGoSiT729OkFiCKFwykSS9/SNpUeOOBR4e/qqHKPY+X456AL7XXm1g7ELlzJfyUNeGVaMy9Dfoq
sc3XLO4hckeGUW+ckA4TLDQnpcrrR8RBEQ4HpIvQ79nYCQhWe2QsZ9hRO5MsojKtWOLTfsru22X/
95c2Aj97xTSCWbQoX9MlshmQpqciT7R+7shbIZ+771kaXk1h+PrzYQJ56nVnNRb6z5m8urdTkR3h
O30DkZaO8dKz696XoIzHQn/pvgGKy+1+qEWDWpsKdc2Ag/QpMUnivYj0rutpQwLithEAV1GLnJu/
1ZSKG1hr0X3M78taXkB8nH6IxnDZ05Y2DguPrXoHbWbXgNX5YI4TwtzYB5iylSzR+dKRB6eCRuLG
T1cKgHpGxVuPSJUH+ZBIvkEjcfEXMzSZ4amlGnKeGOPTqLLYvqRbmNz0IEeP6kindcYuxFdMJZ7H
yfOok3m0b2iGH1jC5Q08c/B/AJt/bBKPPDo6CgMaZe77cUVMP8IdlrmBys/DqYJrOIF/CuEoFgnc
WuHF+VXkBzQnTgpYqk6VuL8qtC9845JGLNtny8ZaQMe3LV4p8ud90ZkBon0Rsx+BfXa2A6oUq/3R
vb41jcuEvI/LGg4b1bLYJfkVlVqQDsZid+tya2yI88saLRxC+96mUPW3mtZoISlLrJd4ZgsV1laZ
1afZlNJU3WsaS9CSjhKa5z0bQqh930QoPoE2w+ENLOEL0u08e5C3fqxhACf9zU8QMeTnRZcJtzeW
D5mur7Ux3BP9dwit5MvuXZqxYBK+FgzWkp+jbZYkOSLCYweIg9awvJmdpYTU7dtDxDZiOucTsDnY
n02qCicJdNFWYsj83Hm+PmmKiLp17lKkaFvzMiorK6oggB7uK6ErAVyhzYwMGYNwqWEodtPaeNwN
5MEQHY3YODo2GqVE859n21J9omnl+ZItSD23qWDzKUp2ekkqLyj36P1GUeOUj1N1o4RnBVvhmJE1
0eghdBacxc69GqLSJnbhYuXC2j+qFUbGm78VkfJik2H7r5G3CUM8U4xt1Y/gBOJwT4rDTEp9BKbL
UmMBLjdpyzq2QLr35eLIopPT8I7eSN7eqUY42F8MtRtkV9LeqLkW9jAMn1UlicvO/+XyoDrzd6cp
FpAizhfJBKhPUvWuJ9P894Gi2WSfBuuBk3ax5f8F2tjRBaaHfmNYgr1qPKxz+IfQM9eQvaJYZLDh
cVSo3sPLuhUadRjV08YXBoU8ri5DGG+PdABTa+zBL5EM1WrAuCGWqP81iqSckaspUymImQKJRySS
JJQcrINAbvRkb417E08YHCc7OPOO4/Syxgjam28B4Lsf8m2X7bhEOmsf0JckCrYY98Ao5gqJ6iU4
s6NzPSSQzIRTKf09lKRrDi5i3EPbM4ue/7hrghSx8Sq/XISwyBP9oWDTkBE1yccRlAfGpdMondVG
h31Cs5LOeyRl4x76Ky2b+h9fsT+hZSY4ZTkh/tEFkFPz/tQC4zPte9hcBLcdyzpZFw9CpvEaSE89
9wtiqUI0ahE+qwx7QkHrpsUogIbSjXVInaG1f9IcK8aXNZUN/kHVwVRhyrZDVf2bU+Qjzrp+cRIL
97n2vMJSZQZsjA9FMnIhySOz6hdOY3nmGRWYbjyW/fufuMgs0JQlKM3oS7iYVmr6prZUce+5tdTJ
Lfl94ycHauOB/CyPjNOj2LuiLG4k+J64ZgEK6FJx01K00U3nYWKihEIaJSQUD6rAeUVXQ2yZEylH
uH43kyp/L5prc1knbt0C4jCXWQlZqUf6ySVs6nIGGuutVTawrGWVMUXoR2qqoU6HtcoZ/67eJCqI
qiNTytcDtzXVcpUfTME3efPPwxqwDQrpWOs3y4/7hiPXCxBg1URJN4ZP8Kd13HqVJrYhqRn0o7Nw
EjKmBnMD6aNrJ39VmwVWW3hi+kL6S//zFHMNB+GBU+WwA+29DziFWO3cKgGaVeQ7fn/skW2UxCkW
I2bcUDVn64/L1TwWgwLWDfEKkBIsczzmjBOi0rSauvg8x7hcTG5vFlHQTY/yXFeGG7cg6WEgeJd3
IZ8vwD9Zr6aP1FSdPY9ffu0i+ONb1jgfbZFd/iHNOfzCOJsO540p/CVWqtnfC54d//zeZsKOxDR2
X7RyqFTZEqMTt3ak8BT2jn3v59Tm6bhYvExl7ReZaOVru2/kE/DzvbXkwfdCS5EctmFNhIXdWQvS
IGJMbyby5Av1Gb26sFXqWIoRemzJUJRD3GauOxQADGiziceHzyhncxbev39IwW2vcAGBs9oi+VAd
g94SMqiRPbpaWzwdpvb/Rq6E22v+IqtplZlQR6NasRouIqc/xUWeVC5AolAQQjs5S5n8jUTPqVNz
/vhEGDLUrF+xqp+2qQsr9ohjkqcLqF58NydFIv4Z5DbqTiy8LSPymeJdIRxmXeaUSMHP5Wg5yUmv
PL4z2/40m4Xu9heRY4GUYNApNDqYJrBJ956wuAdit2ivwMv/k2t+KDaFunw/ghdnxAmugXecr2oU
AxTMXeS+7McYdc8qTw97v3WtpTzJIpZKWSllz2Tc03oS2DWFLS3cR2keRX5DGxYAWKRHZgkwXD++
syPQKPksIwhzFEfOK0t+j3nat4Ybj52DZcDSmlL4d4sHXk7rHFx/nin4JbleROdGbJ6AVAg6sPL4
R6HqUS2jzZ2d5GnTTFmBqq/zJnorDyX1GAGE2kwSVqALefL90f0qm40SW2qrJZGSmIzpOhec+f8c
/gbql6CZeH2NMtzKF7aQZ3LMsS8WRZxd3Q9a6ZmKXkrg1aIZjQ5c/aaer56p1+t6KQjC1K1B9AI6
wWDCxR2U2QxBzWHLMhIFM1bIH11480a38H+eqeRSYeEtCrPL+oo5gxC6gY0Z2Ti0bkmxAc+YXDj9
8ryUXLlRW/IohAEHCArkSUD4cMOmcLeXtSkBqtrnDU5dE2omRMAU4J0u+ywVJbZtbyEBIntoYdjg
Y9T/qMbFMuMdeQj69fE1yjfJt91PCs6XGCTyT7ihYJzOhbMaaOuLCWtTsynrZTdd60HM7Pyd0RlT
T85gbjr2hiBdstomTPJNoDruTwe81NkB0l16bHPyNFgjYHCATFoSXZ/O4hqhGOKhlQVArPqZxUUL
Ep76y9xGjzxXyRt1ZC7b5dzN8CU+/K0R7l9QDmAGrpgve+N9lKvNAVpwO5mNAOzZXH7gvJjnuK8A
lRQovsyJ38jJAgcdQSboLk+gUUnrXXJRB0+tAmCy6fl00ptbGwRAJF0VnSqn28TPGvSeS4d4Qas2
N4ja6N3zUh6d7k/2AnmKC14eFvjI77jYQ6Y/lwvl5rP+XqS2AtrD0I4AVZeGIOVfdX2EEMiclqFx
P4omz71E9UbQ72iGij3aB8hipdoc9Sw9XHKUqSTheWT54SPfD2+CDZYT/4ydqnC3hGZWBinb8+qj
o7YgpPYHeXFQJOgtHkKzXxPPqFPt6POVUNcGIJuSzezOzBVdWOyd7TgYxKlYr4P2/MIXdt24zBsq
3GREsXcunHVi/A6gciefkoKhxzrhe+7SCBMT/mziYSDgStudA8dQRFK5izKbAVagfX4pPD6e0DRa
5UjiW3S1yVmgXOPcZOy3evz50I6Nx36HHBmlg/KacfSbyvLcuFqNwSfTzW6IISncrpHDR5u7bDVo
9PJJNvP+ivCqReu2CS1q9bffWmAMEJpS9Fe55fwVRlZT0KJ8gSWU3+a4oxhQie26QhVgarbZ+CQd
0DfJfoc9AJYrO0gKNixQjZHy2Wg3yg6NyPW4nYdW8aBeH7ZQiH4CKFVmzqFK26oqdsHz9UhGQzIK
D9pV/3AA9zlrpbWd4bdZCtvSPY+f+usD1iKAV/kOFy/U1jI29XI2EwLHKEdD7VF5gRrGLTOm0bnw
bDbSg9M57SoDimWr76LUMAPESwgARgYKUH6zfvnxgw40nbn/je3l+hL3eOPs0YPrBBjyP0na/63B
sY3mcB4vuEKycNFvpKEzi/B+th8NQl+X/XvXoNQ1UfAbqE9xZoKSGrXJEG6s7XoXScAlgIRY01ca
YIbcEmzr817iq54x1UgBhbEQIkMyeofuf6mVqmIlsYJFFIhV3uSEnv41Oozt85sFs4cOfhqNiVg3
uQh7XK49Yr9egAuwQvWgIBw0DID0OcinRFs6MEcbqb5gD1S7g2+AyLIEQ+m8pg96Qa82yT8PqsTB
CiZ5R702HgtZaTcE+D+coIbE3AKYyX1ZyiuxeGhFaL5+tZhIro6Xwdt0sEPrLqqjZn5h8GU6vHme
H07Mh17K7ipdUOxjEnRIuSG9oiRBFkCkSlNSD7OVo5Fc29OebAz0rEeBYj12ZnC6hUub6ER5eEI0
Ak4oCMYYqeVJxeyenV2J+hIIuwJSYaXwRdhLqtt68ED6M1euw1JKUkYMAyBaH9U00xH2NnJ9ZQk+
544OEY6VifLO+62LvRH+6rLwNeWGRPc+63J2F9Tl+nlzmSjRjy6cCLbIL5BkMgNU9gtPi5MvI54S
m/hjfD/k/NJcp1jWaowpvx2ojvPURz6mVvzxmtyGkNFKy/leX3DQfVmHiFvlQCMIs817PaGCemOP
n+exUrio8D6XFvM7XIn4OzOBv0ZvOSI+744ZqVbsm3Ok2BvMgFNMMWhq44fEOqcI+3LpucP2Ow1U
H0cDe53qtB+4tV6zVBbQMAeC0cr13KeUB4tA/s5SbkJJlV83R0VQdqYVovrPOhsXscfoa+YZGH4L
2CR96OlSLVwFJsa5sRW3Yiur4mHBiywln6YdxdUoYFfDV6lBXWAvM2YPR7KyuvCBcVEKMqHdjsMC
wsaQfCeyLe1ZpbhxjCBJP8oelB5uJh3g3+nYrxm5ixx6swLUAKGiG61xq/xMcBTXYQYiOXGjVxpr
BZDN/yW1AGeyVykyB5gQmQnJISiZZXX4LlEY9vF1NaYj3f26tHZ5zoVT/2Fo7Ybpcx/MxUhwBJ5x
9RffoFC+zmK4omy5MNRMnjcDgmSpye0oELOfXP82XkhBBWQ7a2pNKK2UKFEMiHO+/hj4XCdSHyrj
aPKCUvw/3Qvetr3t7RUtIRkX3hy9sD4JeihoiyPX2U9pcGPVA6HquvqcvzFxZj6ZPXNA7PbkhqKw
vBPEbS+lOOM1i4RSyuG9B5RHsIGyW9aSwyBW5RarNiPFSb0g9b57bu0mTYe2nzCtQVusO36UdyxI
CL27O9HcLUT+FJ3JICxQckz7oRnHF4QoUNybdPFbjNHMmFVxSvd9WtrrwGH8JqkY/T/NjKfYbuTu
Vkb7pWr8e8Vlmd5/+whbrNlcQw+9WneLSu4wA/eyCwJYrZj1Q9fA9Ll5hK7BvOW+SnQcIbfQynRC
QYazvGp48Ud5S9FMnUYHm0ywdfkRlvLIwcJ64W4N4vRx0g6jMHQaHvVQId7YRsy/EzuiX3VYoQBE
3A5i4pPUwJUhoTFHw73YyY082HL8c6OqvBmYIRXd1I30wI2PaGSvPnYHl5SIIlbwjhwwuDSZvjU1
Q7wLKn70L3DYxFu6fGxLkAQPoyIjTLPG2s0Izc7hxzutKbXsp67KWL1+4zj79b/X9gs6fXbiIPeU
mLe5aXl2ZRK0zSO+sqJjFdGYRWHpSYFW45JpNsHbTu4wNMktg+LnNeR9QVBPBJxLHihCEc9hcUzq
VzvuLxwfXxyMgrezLbFx+umfrtVJv/BROz3c2Aq2nHCRCQYm4u4emp3p4+oQU4c3kDHXuhhZPZIm
tfAgKWQe7As2rabSXgv5sk8RPdeqxnYv8D8cRIST4PFc6aSTk/bkJo2a4d825Pw4x5Kx/snQKQi7
sUrO6vBL+1H9px8CMf0bcX+ZI6QWWSNz6ZMqOxW+BCplf6PJ5NBu5dtM83lBLhZ8tkMFhTGfhmEa
52x1f7Kh71+qGTE5qhD704Xcb5NwkI6pIcInxoze3xfGbpIHhFS3eSKtQQ6EVjyWGDRHzpk26Zhc
PB/48rH/obs3nrUgBzaBaWJgaDBSsXeS/pJvP+wJkx0xFmoD49NLClaM5e4wu7ii68Md1DSDX0D9
IEBTKM0R+Tz3cihkp7/NZHi2SndcbuGqvH8rg6YlfhNb7XtpK4LOzTArkY8/rD5t3bu5cJaTGNYu
b5CAkTQpG9sTnvHp2zzlywwc4AZhqFsSghc471GdkIKwkNu3fJgNhCb2NcVfV4j2ZU5BPrY6OzCx
RyRTHsxwNuryHLxLVEqWY0GkqcfuL73C5OOZXRi1TC7ku8/rD7iJiZlLqrf8sa8ePYdysDSdt5zO
2KYTjfImoYGcCekfPM8DhlYx7XNwqtA8FWZH9K6DMF4jNgiT5gHebQDH9E9zndMs1d++QqUKtraS
X0oe0qdqDRyE79dY+2KoMBE6tJu6hhFrJihL4boczZb6h/YsJvv0rZ+KkjW2b+tHuTOIUNmJPciT
hBhEo+M382+7Fzqfz9xJbu/pWofUig4D2kMemKqjmEk7s4kD0kZlz938wHRCE2CfQeWbSn7UlaxC
QLz8IpdUadjC5QmT27t56sylVbfMvj44FEuuiM012lttxZ5tbWcAanfFovgZZppXS9WpsVfm/LXK
bocfoHGUFHpLb1ig0N0iupMP5cdPFjtI/uAORSmVQgUbzcVpvHUbAEC41FYR8FlmBVm0PumO5IRP
V6MnxdeXjZMT9WA5cDNe9943flL3HzdM+Q6A28IMYmTei5YD15vo7F8a/88AtGvnwbDhb1AMqHfm
Z2BNdcYBnEWO/UFEQzcaagkoKMxagNtgN2mpaOBEWxIgzXmD8/e/M9IcAF6eZDRH0YeQdBpX+6Dj
b4cwsjXU/wV0Q5sGbOgDB0kNZ0wqK2OiuaSeptPHZyY6vZq6jcZGXRRBhaENvU0Kwu4RGvxzQqeD
B8W7BXU/kR3XF4+ZdAxLKQdRwuPZa9UXzk7Rx+JLqX4YGXYXJBdiA020gI8+1haQFj+aFu2OH+9H
6BuQao9COIqTDDfNP4TuZTWzKtZF7fLmUfwJfbTMXCLGze5DR5vUAcaMDQMU17hsYVxtk6YatDZl
CJzMxrAw38EmfluszNzshmytt/NlA0Kiz6UXlbgKX6GBzYpEVaYY4iKWKaHyMUEjcfDCabCzj3u2
EkWAsWqvxdUAqSVRF5PhYfpXPhURPUHM+bcXAh2Krluuw6/fPA/LC6Wc6Rhx+yuGdY5B8vPrYimr
qZWJea3Usb31YFP02vwntEbBnCAVxSa3i1I80TpEFIH9FzsnySZ5VKFl2jg/gKcEPGfnHTTNgQ4G
+Y8MTVR7uOX9IsEh+qwy3B7f7OWP1A+IZje+dW3Cwp4Xs6XKrfpCpaBNtGJYIXwR2gIA49KMyRxE
hMEF/RdZSBp8ixOqzi98JCAxVVMCIfQL1dGVQk+lTuoY+95wL+ew1lWi5hRyyCfEoi2ltCNHyBex
ttqffoDSjVQ2g+j3yOy7JL1uVueD6gCI+G4RzdMGZ2kOs8HHWXHbPb59zwij7Y4OgwIvulqphRmR
bN9PleE24RGIEahJAOwJGx4OImiYesEHEKDLInDH2GYwIA/iCcXbRFhpaSlVALinn+eByCLSWprv
qrWmJfd4/FcN4cZSifSzGKxrwbVNNaUNJUwzF+qmTuYPJFM5ZySqEOeX+a3UDwLspuFE7M4RHwCK
BMFiiPGuvkHALSSu3QOrtzKe4r5mfiyJVA1+eiEGQIwmw5NU9CByMnyXd5Ye38acaZru0TdYNC2D
bx19EyM3iigMBDG1APF59alXI/I8N0fffl0a7Fm+Q4YR7MPwdcaO6mHPhFwaPdw0RKacMvQU7hiV
sil4RamJlBzVEEnxN5hmeh8V5O+HQGVqs1j8rYBehScEECXC2sf9UpAVcVdYgZIThGTiac2kG2Eq
x18Kdr6a2nSOakF3q7rqHwf5FtqS2/b0gtxUY5r4yWTZfDoJIlyDURfIhnnoHa/zi3QkSYLc9QYT
p8eOywEbw+aNBj2WxdJFbO5iy2hVz+HLEQFrf3YOJSADSiubteBNZnHIIR/+t/i6jPDUUMjEbKmf
u/XqZacfXujSO31HZaCA9wfjoxZP8NqQvSMMoo8k2Orw3F4MjEKKL2QQV7ZNiXKrM4AQGl6+Y1+Y
aGfxzT8anSz1Gakof7M1ABuWQ6ocDXiXXECKepwjsJdLbOWDO2FddCDBvMshnXJ1ybikMBRiXcEq
5vpDrYziJixiBxGxhKvGLMNWfCVoKWB0o+QKseDOOAVPdR74bos6On8dxj2P7nFsjsyaNbLYl9ff
+iSf5lJ3mhzDA/HrjanNiG/gHPQFZlr3dvNuYPacCy2XyjgQzL35JojoBnRgbnenUE1UzQxlykcd
Qw3s0yw5suQQmL0CjgKUA5c/QWH4KTxOX3REaqRWB/PcBe53DXOrqSTXbMuK5S43uBoggk1931Gz
KBEEIoVSs0LJsfFDDMKyxGZV+KA6YRxoZIzW8t76GqX/z9NtuhAyMihYLRV3lmkA3PfwTQbwd1aS
EOSWaqxQEeC8M40xIuYDwbHvm8X+ch7h7+NGwemQH7oAKA2gXelcJ21z2hoGE3kqchIrnSlG4Im1
kCg0U1U4BXVrv6JP6iY0lOGNaauoblAGcjI7s8eJ78DZswaT0QA9a+o0qLdigzym1rYRXQfAAxSQ
sOBNwuVeAmSbQH8Izi1q+49bKNrEugVmzU13ZizKeU8G1S/XItfEcKdo/v1I6ZWVrUSLixuO6Aje
oyhAiFbCdQUzqbsD2yvKjIF57uugLqBUqDmFLE2JIDEaO+0rwbqT1jJ5bWWj7BWGkAKcFRCNLYXj
Cek7s9VPFV7IoHXQ2aIRJiJMhO4zIkxmwDtm4mUiUOrmih5egoDK6Ua9WOTPVevm3heGSJoY7Ftw
MFe4//pfECYalEIeO3V9Bnv/JT1fLToslbrnnTRGgov9i6a9G3aZ4vaVhutdIVcCb78f921y4nBf
Ux6Kd4+ArM3DxA4sUBpFuHpR9fGWr0mfW65cnZjtpA4BcPjCowpdO5i/RFnooYPCwP7W29rSnrWc
C1rnOVkB6LTclzjqN9pQcW4ogzQqRDNBRmrkAFsvjRx+7J/TklSU5FciGFJOLf/VeMH5Lq04LmDd
9VnGJH1ePqH5Rckdhr7DyLGBY0ZYcfEPMpoUw3dPfZG90taMaUAlm6v6cwBJpjB53A6nzCypkeyU
tBowAtQ1CqON8Kc4MG0H4Jfs+rlhiKCS5cyQwAk2NpaoTsGG3jajucKMCTubrVRS4DcsrCgkYr6u
GjeVuWwnOPCx2OgpNqUkXAprf6W4iyo7ZBMufpGXRQtJ2FoDtDDnQeYeRduTgemLdnj3EvOyIumn
zt2XbmjSpPOXq19/5nL2zBTeQ1501ZR7qkvyYq7kBjwAlsbeIdqGkfLDfZojgjyTT4zcE0n1xpvf
p9pLTnFX5v76I+dmrbZyyKVgIPrIiYAqyVJa6LkHSO2+BdGFpieeG+g9THbT3gpyVo2QFMPqXbMN
JOHKay3YdPLA8Ua6xJZc+p+fkIwMqFLdnZ3X+g4hNHpkMh5jNCoIBd9BCXj104S1v+giL6arzLK7
JHaCtUZCdxDnJwGA2EEqpCA2O7b7Mvi0iZist3FBbXZrAaN6UvyCFWLFRFrem8Aw58rrENMBcVwf
9/OBVSliKkSZ52tB4X7mZyoiqP52xDBniOs7syw99xQss+Q9G5VAj/LkKLxQ6LzlUrse5Z4/ANEc
b02XSJS7Zl4flKnEignd8m4MsCcDFhgfWXilvKykhh39/pB62o6NjuFuggBQXrWaryGRe1JXQBmo
uoJJHgL79/sMujZAzPOH2e2eGoqrXjG9Si9H3qI8HgdrdQxI2q23gdrq7T8zsiy1pna55flUn2lP
q2WduMWMZhQzRexMJuFmVJJPTzDNr5LEUhjp5rDt4vLyRwe2Jsfdcqt7B0Ro6fq8COpOVjqj4uPw
8Rv1TrO2KrUtSpM5Dza8j6y0oB6gAD1AR3UnUzxAYh+uf97EeiNcq4MbbZzvNxapAq0b2saKbdMr
e+Wgs536EaBBG1+0VcIBs6OAOJ+gEPDFdNT63MLE7ksBeI/st71GR+N+yS47DgdVVVGk310oS8l2
dM4E9dQVnWWOopLqK+RwRBjWgFnssIisG0sOLhUbVTmlP/LeQ4VEPUoc8X7evOTHAs27H/dfoFTg
5UX2tSflxqASwph1OZ2apE+fSZ5SfFNhGJypr54GCX5sSFLegmsfsIQJnIQywSsWA2zoB/DX2hY6
vbWaEcDeNscLacNrogF9sJ9yvgiGE8u+FBLdxsynen/dC9ybdL1o26ysswDmOD1p64b7BALlvdB7
nTM5Qzikw5U4zMRwzySclReWTcyix4BYRDNcTaiGHl4cAhUthGq9gJR3KpclDV8XQkiG2r9qGeqF
b2iBuY8+6XbxsSPF8c500RfxFmnd4vpXfq7o8p7i9/wNvywAv7u9eAuaOmk/ng4VvWyUXzewgoIx
Nk4eP1salr+X5ttnKN08/AQE02g5U37zc8z3KpMfexqz9RsdQsTvnmPJ+tK7hrrrcxpaC5huIWRJ
qqXfV+3IZkR0ieGXeEfrwfrKZXWjjWd7rAdPZqsZoVeWMt8g/aZfkXgsHf/BJ4jMzuZOm7aJOgfs
f5IOWC+IgWrkLl4J6h4eQN67ngC8uNOW4A/zZxOtmjBa8V4ByGvAFNaivapf3PbPe5PosoqTAILj
dL6vPcpxjeahP0BT2ltNpWqJXAIn8VjAj7GJlvmSsHgfx+Ao3JnIvyDLVb2vLBySeq3sj18yUQCM
NAr7W05svRRy+3cT+44wP8gPJD5syvtO14nh0Pb7w7RJ3SAJsG0qD9OS1x7EQLtvdsTIz1nB+aYl
iB22kiezwQpgZt5BNBP4RKetlYdmfdS8G6F8WnhA6p+kasqLGmGCRCjfyy0t6bjFOYYzx3/Emnol
/lKN6UVSGMngM701rw5eRMc8a3HbWC6JA01Mb+nI2cpYEGJmPRVwV5XrxWwkH7kKEZ3EzJOkc4YQ
BeD3K5cKeQqinf/W0uYY7iZ5UPrEI4fW/7XP2sny5d1lKyBecGXBPgqy+4TXk9NVQdwgjb5+VZxm
ZZYJAe4cUROhRfEMgL1VOQT40kLLg5iBQLrkpKghE6VAcz6C17JkqkUCRKtQVyL09xNTLpTjAswV
e0EI4jhNJkBVg2qYq0GKPIVRmQUvmZGbt0UBAQbDV8AH/nUfo9o3A9ynO7zymicr15NWZz9VgM31
mT5ZhiOVUtIb3GG+1skvCCgojnbpFhAv4FuwbJm5IDhha1LuNRB4VRTAD53wdcwMLKtasN3vhK6i
k07b7FguSim4sB6GwkxG329pSCIx2Nk41amZjOXuSr7pi2h1RnQMhCzTfMBYeRQRZ/0AdtgcLa5r
WOT0a9+OlEqgsbsSjvDenNJ0jOb+iKaI/ALUVpzA0epi+k65588MSmKhRJ8LmzvJbrnqIhHaD/nY
+lSn3DFRqzajYWsy4whewMSNZHw88mRpv9bAMiTkZXpNwqlgoBbuLGblJwSodXbR0vnPi7x+7tCe
UNfVUo+NhhgF5cv1ni6Cls2DyM33hFXt6ndK04jtNetVrVttbRyo9lstJxW6GUgHXIAYSDJHpoGJ
vS1ZBvKshdUNe/Ui6XQ8e4fKZy3hDbJo0P+F0ULiP2CjeNnoJ/yafE8lO1RtXYR7WsXpss5e3gxp
lSqakSOQwzqtuBO9uFsIY0RCzIJtbsIz2XiM/Z5bYkau7De/4oLeY8ePaSa/kq1yRAnmONtVy1zB
JmECQ+OFT+oNAm8BgiyCo70oXS1KzmA25/7ziLFrR62qSJH4seyJjcG1O6g28TTQhitb9Ftp9Xja
YBvXoO4v1azD+pI25/5ZetikTOw5fVe4cPhcSDiL06Uo8EUBm2NpNx/bNC+FF5PByhmJnEfZgr9i
6LUdBAWYD7x6H1zz7KBK668qwgtzyT+zN3/eqdGB5WDHU4mE6akzUyUg1Ug3WWFr/BYH4FRSC+tl
6lrN4WE+YWz2ji5kD1n80jMVCSBMBfHriKLyy0OwaMJzJL53pqES8a/Syus4ZobOWr7rdfDkezVF
RaztpX2hH+rJRwOdYXyX1/SXFSVO9VgaEXSLpmpr5wMgdrLX0QL9uqV2okyXeU3F8CbFJ6kG60Hv
hfuqfjxpFObsd8rnNg3WgviMxXs3SbG8XWe2Yz1/HkNQEr9qrVf1WVxb/O2Ioy9UH4RQFXEZfPf1
R/zTewys0CM/CXtxI0dx9Jdwc/y7EovgeLQeRMlrMnJ0eDkhZTaXU8aBFZ4APS+7DHJGCTuBq3j9
lGZTKucVA0TrewqR6KinMOHNlCKRSEdizg76bxoM2J9kYK3j1RiKtZpjwpDZ2e+NwQULM+N2z752
tfeUug+frjJzgwYXDM4JsEXKkSSHmVddp28iN5ACTxUvMfPipu6cuNLigc4EXB+C+M2UEDi2FShh
WFlfuRXmBsL67lsebwefds4KQ26BiV+uUYBC07t0nxocfcSezDKxdCXhdVv4mdWEqf/3SvQ+GDhv
E36ccZ/DrhSpFMzzz1KCatgV+UkxdRXqu/ssaLWO5kNGqW5vTJ0qplmYuycfo1FsVVs39LacHSlj
xGSkm3GsuePA0GNzopf59uaS6m2SJywwiZV+hBP6ofjU2GbNceSOmd/P87FAb6G2G4Luesyr9Mhe
eTvskGAfl4tHkO71x92gpGzBUH6tR+Es0gPRbooSeS5U2UP+jaH9rMMQsoSyWXmCTNc8/vKH9OVj
Z130FvwCIIHIqSp1Dtk0olZF67kPbub9BDRONSKgVkGM5ntkAweiaSLEBEMuAa0Q2akOyhkdSfrR
z+BW5qQ9XyJ1QD1bUgdnKG8eAbNx3y5ULtraOf36eEqeyY0j/lvGK1Q53BHhjCz1ov1cpRAazxnZ
IW8RP+AmU6v+gVr1KiZ5TdpxbPZnzpcGDJ9uXPSymy7sjeAWyDT9l+m0jysstt5PQ+2uWDniPZ7P
4KlYXP2fvk0DbAITz80jw/ViwDVxQzfcijVVlE5PuZUyncgoG8z1e95N2/W9nvYusBWP1Bl3X7S6
OrHfYT+XVkkDqY6jYwDx2EYe4VZ8OpGT6bY6vBYrBbW6unRkPe6wPxvummQfw4Ve/iQ2CWiGjm2M
STbDbpIDvdNxUMAj+UvosIQuktj2Dn/hBrGIlipe0IIstp6kyjsQqhVmpYr4wl9m5yvEA4OKz91r
AxwK7kVi4OFoUpHSE0VSgj/e1P+8Eipdv6L4Mp2QAT60h7OjcMF+qoqVeUPNkdUG8Z8y8fZOJ/gG
Oko9/ihm2CqFh8n9RQpEefe0c6AKaGkRwJqfOVKWSLGw7mvmiuV3MrY1Sru/Atzgib4KJtyHO0no
2BfC1vqMg0T+2Df5Hi3odCu0KqtQKNIrLE3lwWboe7lwbquWEhao01u3WmxthjcCfUnzbM2C0fkN
6GIV2f6QF2EsquyzIdV7wqTjIz+smTcchkigm3zGWeoEcT7ObUAaHF4JClsiBBxMIFyt8vdE9wfC
PTVKSXBwwsN3CRAb91oXSTFvAU5pe4SzvebcY8ob2Nk8PsyDL8gMYdwwEAPMEp13dE2/2/qd4nN9
8nNEqJMbvUNzADtQI9WjVkbkpVSJawAzaricuZkSrKEuTx1v1AiJctgtbUbRyENhNIlNNwXosIxt
GAwZBbzFxdrhp6odz+LHPbMEQ0MBe/B7Y8JzMOcSS+h9H3c6zX3/kvcFdiiYvPeuYsxoNa/KG33x
sc9YJsUO9h41ifpZvkht5pH0ezm/F2z0ZSprkbVspMjXhCN7dZeGU9brk9CYrHOByONRpXXrEiZ3
RWo2NKpl/xi6qGzQ/mIgSOpe37m2//hNH29SSi2qS0y2sR+emhYVF2RhWPFF/BuhTPxmZCkSzffO
kGUc8e62yru24GnB277r5z5ej6Zq874BsUBkYuT/aY/cTvtlzRq/r1b9h20OySDulpfcRGkQ0NWy
uF2HaV1MyE63zCBSqFFFaIKyw3NEN3CbX2St3QTYyuSP15VCmw3BGqlsEBOB4lHgWmfukIFTatNJ
nl0kVg1wAZi3QfLLnUzwc1cV9H80l+5lnNulFhnJHKxQyj/S6qegp/flsJtatmFFMTvU32yP87dt
j0Ev0DDJhsM2e4t6bHTcwCd3sCkjQigXJKbRxc5maZZKu8ZFOW8soEnik3D8l60KNyo7aIcf/9Tx
fzt975keClczbE12p/4sT7Ang0neJ3ObZg4oP8nk404B1bJvAyTCdwNOffgbi71KkBXEr8glWBwB
+M59cYRXoH/EMHK82PtTq0As7UIeG+Bs5swdRrv7lQmXdC5vM5c5tz1v7qaZELE3hzAnFxI3B4zn
Yf60Hjk/ASpwANDfzMRioGbRdGnWNahejzUt3fMD2RaJ+PtrUxXR3rUP2vVwziLgf7mkKLkA0uux
GyVMeawbzZajaQ9C9CQ8UGEuT92UJyC7gCK54XZOxdYLC/a1QQqBOsYMNStbjvpaIQJipqRtszZm
a5XNKCYpNgVHw64d4es1cW7gCh8nRpiu0s8t8/S0njGOC6NIO8fX2fX158cEbq/iVckn3cVhydoo
/ZfK0sWoyMZXeaGh6Un5GXzoyO0YFrg351pmI/dT6Fvmj3rZsi1WQlAEWWXvuUDJ5eu8yBVft8je
qopU+f2BXP5c+UPddOSrqQ6eYQh/lQTNsmLnmUYXvX9/XzliuATFv8mQ4pwoCYlCz6JXaVGn7D6W
ettObDSwiEPPTZ+Y2ecwn4Dpq1nRMLyYyHRqK6dTHnQKBPLP12U2YBD2IjA3z0R/m1RU3Xbbo8X6
IO98O6ndZFu6dx4a1UA8hSX25udRFMouYeLbMGn68/pWmy6ITC/Mou1U9eP5f5TLiGClzijQxGjY
KGR0sP5UZY0U/KXQEWQg4j4VQR+fpy8ow6fM3d/OgnBaiR0S0yi88LeJa8atOptDwed9bQqgSGT5
Bi47sxeWHIZFA38Yx6KnZabyvve6ydq+a0COeC6455+lirQ3FGCpL1CRGJiK8KSmuJ3fUujQ8hCz
ymhCMZwLDDMa0L/jBrUYLDsfUC5VY7c18rqvenlnTbOb+BxPpVMwT4TX9GJeYSt0tjgxadTlqzay
masCTuRDozH3lO41uY+ewr0m5hZFLTQBRT59i1txA7J+5WQ16BYTxMjomw2/krwTivvIn0l+xYPp
BCcul20pYf6CBzaNr4eaDID+K+HgemFio0U1NLuAr7w9RScpgCr7nW98tOvp6BKfjI1CUBGD0PKy
ZyNvI5L+ZrG2fqLwGSNNpn+VqdFizPBCAgr7cTgVtV3Goid1Bfd3ZMoTbB9LC/n5rplBW2PMCbk+
7pwnrj48+d/jNgU9OLaa1abHn6oJ9ngNlFXLzogo1m6Q7/nEwnALQPyvZtRzvoubuvkqnCjaaRsy
qcLQAXcczhb3hdH6EuDfelemc6+W015diCYHzSGrsYFtftgw5fbIXT7pe3twg9xhHCx8fAZb7XK5
lBxuBnltY8WX7mKEpKKxDY0PSk6FIsq+ZEK46He7h7nUGHOfAlLtPbYzJwRKZy16WjglVmGrYoJw
NotzpTrQPDAGOuKWST1rfBB2vlgkpM06qSAUlRvBULGIJytWQWczMC5SFibtIDfbxw4BpR/+H+up
Odc94owe9JZLs6+EXmWz9bbYJtIh1VeCrvNjapmzP4GmSL0NLPrrwQQGfOUYfs1zVpTWqiEeX6dW
BtAg+9ftT8yq/FyZA9eE6//cph0Xj9kbiAu1mxmopjjQdpTcuv5dV1D15t1vE9mH9aLp+FH258b4
fVcXHMqQhGFwC73FRIeQym8V9IWqZyjcZizCPiHJu0iPt2MkjO1J4lLLpqcieJUYqufFJkahDWOa
p5hu3K/oLQQon4YEFdEwRKcBvss/XQLu1yOPwFyoa5KcqWFCPZKPWS415nXTzFiAsGdLHURb4M9P
GwHd4fRM1i1XfF+5/seRUxsnSAZIhSDi6KcYdCVXL6wD2iqzNcKDYJBDVTaSte7cS4r0Ag6KTsgR
SQj8bJQa6CVt6X7+NxdRwUGXpL8mwrP4sZGl0wke5EE3vaSLQ7xudBYECprwrjz1cAsy272xXbNh
Tjwji0xVIqaXMEvn1l68de8nOyRsNKgnV65tmrkQIJRClgG3kG8NK8qNIWUpiJjD7jE8yDYTMhp8
t7PeXRo7rL2OX7D+i1XGlH3AgIzhvA7WNbBKlwKVwlwHe9hrJQgbpyjgScYoSYsZfdMAqEDtFpdb
Ul37P89aIaKvlb7fsFCGBPHpwytkC60/pIjknCHx+FoVzNVc+wFqmWNL9cfBqUpgnd4Vexey0Lbt
SOM/jOdWuUdy4VuJ6TpdeD0TNet5B70Ot1y8wh5H/oiegIEzExtxun1zhEY61ZGhVLvVTd2ql9tH
I+r8/OOfNnSYXRSOb+zMTgRPp/UmS0wt0ERIY3B6RKsT8hXVKvzyWwZxC6a/82GFKPapmOxXWGpZ
JLlv7mcfbE310m9romO3qBF1V0BCX1/VL+iPLmJRlppyTXPobpsBxCFT1Vphif1nFYfP0K5ngG/E
14P/lTVBJCoHfVF45t1KwZPp9Om+0uEfzhAA1r+lH+TKkGYZyrnapZ9bequ4EngM2URJyRWOmQCE
gKpAAuYqDinjzLriR3XwZwUgKtaj3Re4AM3fTMEPwo/jyScbUQM8JkqBh27mz5Y1/wgHiRezaCsR
EXTq60rkkWuwIbV17d//s69Gx7wy6UT3TLCAcogGViDGezJiUNTdAndAH2y3km3ER0XkbOc2iEqa
YfGvL6LqzXHPRGy4tZLXOooUvp9Qi1ZGnS+ceddFc72e0LxfE8HTASyfqi0lXpKT+7nTKRmiMgBD
/Tz2nPnQTWXkuRk4uZmybSWvDt6JmfC9UI1kXCUxOkmVyvbbNJfTTfth0bG/5jq0pWpVlTzj5+fL
YUk3W+h1jnWdiKw0k1jIRpG+tLPvN/ZI2vVbzl7DqDaVzRoLNOh6Q0dSP7ev91larIz7QWykuB8m
8J6Bkoxy56pVHFbpTr+FoaAqL0aptDGMwUex8CnWBUgyQQBTACb3zT8NqkNPNVUhgUiEoV0bLsUO
obHNlgcvQrFsgOTttaExRBD+JWE4Yok1u7ZBepP8xXMxZvMBz0eeRaUEDG1mINq2FrkLXMs5GdV1
KSbx6KHC0QM66BbSM/sdHs/RCEsRuNVY0RVLXNto1e+PQUBTDYsPcerowhMfl26hRDfavzEHGP5u
NKqxW6W5zR3oNXXQX1i2uvung6D+6qK+V8ZeooNJIvNeNhIER7Ioe/GKr45iaKySpkHPLlCuQPgs
sgh63DA/jUblpVlFOLvITel2hJxMv0IMHBM8zqtz+B7eKhqs1tu3OFoZYO5TI9hLjwbL9ezMK4dd
SjJaoDNwqRpbU2vzTW2HYzKKsXc8lWycziq9eyxxzOMkbTTyyO3AcszDyfPDxCS2BuKfR7kz6BnT
pZrfbPr6P32prpHsEdYzpTdgoymc28y44QpAeuaxTnyybCYSW0NILPqeeZ3wrG6dG/7/K2MxCeL5
NbuUfN4J0KenFfYzJeChRxBlhLuV2mf4G656tcIluSt7IjZmxflHzNu4Qz/8Tn90L33Xcz9xtPga
dqUFTzNgna2uiRxHV68QKirLgcdtnJpl8Bbpb+W78pt79xa/FZfnfRcaBe9jpxVdyZIhT704kxyQ
fk5a8qi88jw6yqBEN0Ia/ZvySf/1eNeRqBdFrlIU6iumpbasGCen+nC0qH4YGcwZu0Nb+PFBqF+e
lOZZoj8CPMz5c7xi1dsr1TIvLwqxnsKVMoizIrIXkNJ6PuydVf7ssIKatriIsgJSSt9rXqrMWV04
0ffAxgpItnby9tukrM1MZ1zGSKfg0CW+C9hq2j7h+vVWP/pNg0uyg6KY4O0dSqPV3WvtOVHwXlwu
mRdgwEkTpTWbts4GzOr2ptTIjcLIW1ZWuB32y8g0QruB7NSygkf4MCKgRRLVsBeFcg9LyqCQmWKp
197enwIzlA9UYyQyUsjENlonepvjUgE3jQbEJXbD+Aqbf7mykuAknB7v4PzbzgH7k0/uBeyj2tgW
hYLDXZAGwSiug/uVPX/HT0DbY/WK7ufrTY8C32LPVnFsIOldIcR8E73E0cCKwZ8qiMG/PZWofBpM
hhdryQkielm1ab7R8nUR6HRVE2KNEZjgmSgQt6NGjzYGJIDA7xRaJ+vEoyfWmwJjHueKwx7eQSM4
KxikOdRwrrrU4BlPRjH7qoqi5I56PYD5Wu5RVnB8l/PzE3adQHpXIjXvTWwSipdkrG2nkolqU44e
pvQaRj2aTekeml2w+uN7vitOnuUjKicqGBO+Q84Gz5UOBLxyhf9L1HPQBoJJJ1HiMmVEpU3t+7lW
0JdySzpFBUnImLJQIgXEgh3ABGqJ4zw83UQ+oxCNLaVls5v1Y3k5UpoZVwJHp6qBDk3YIPj17hkq
YzWIUD4nwV5UcLXZ/MHoqTUvSmh6MICw7ZwC92diyzz0pDCoA9vhw6QVBPKIIn5e4arTbUxWeL5x
vKUWGQRw8zVJZXgDeHB8zbIt+lDi50YJNIw7voumCMc1DjrHX8jfibDgjn3TQVhZjvqvo/eDu4Nt
aH/ABxwuMpdClikTx8qkRG22jT5aipUukK2OPB9fOZbj3FYYsv91XfP1YPJG5dcSVAx4B0POnlfV
Oo+tEBKHL2Ci7R3F/3c303osejEc8kXgXlUfrPyPiMj6nU+CU9K1SsstB5Yrgspxe7VGAmpkLZNj
cPjdkI+ep1r5EY39oBd1at9MqbKFIgEDjBGo2xIMEY6i3RDF9rmq9/Ghys+PCPmWyNbatleo+oL7
hlSN1YN4L6+KHj+FLU0XCsBjID0Fk0uLMKTX70Men0ULUxjgPlrM47GsAtOoSJ4EzEblKrjdz+sr
YG9FkhGmLoPdP7ghVyDXpPV7Bg1NjapMOKfrC7B4npDLed/Fdp2ECtvTDxFlhPk/kwr1kD/sG9uM
5P4y2wttzpEVyC1NAAmG6tEtpVUgDRkoXhEnSvUwdxD+kLIUqVyp1AKkA0Bn2Aa1263P8A0HwlgX
dQKAPpmbZIBWjmsT8wNEKxmyEfvHJrLuOj9ycyBDjI65w4CqFgxl8b1LwC0eSMvYF5/MR1WcfkBk
CZImsy4gnqjyWLIOfGeb4kA3/IeRj2sKQJCzYEderwmb9Ljw9pUv41MR6vS3ipfG0zhH0gPzR2Kn
tZ/Dx7vT6x6ebEd5lK5Ik2kVGT4fh1PQTN0e3Vc2+vQNO1bZHO5oooO5pxLO+6G4ImM43YQPbbCo
krTeABjv9qgaQKb2NsmWGHq6qBInTtiaf+65YYP2xkpxjJFpEz6JxKAsZmAVMDFrR91XilGj2pyK
oe5CvIAxQ/SHAPHRHditjn2SY7iCpFjFuJXOZH53vWfDQTty6ah/EBWAvrTjzkYCm/3zx85sKS12
kimK9TBfwrhXoKUMD5aobdcUB3gAeiYW91ChAghgaxvTEpOTMhhQ5hwxLjmz/yii5uDRq0j0X6ZZ
2cQq0+7EFbtbpqiohztbtZxJf8dNfHUf7WJJ4NuoZ3uwFS/HGvXE5OMW/cCWRytGHrrAx9qVE9+c
l6iwXrb8W7jij/5DsxRKjaVkwNkdpyFpqrNjO8gnYrkNzfI/ycrKN+Yz8pYBV3bG6LXJ+YzL3dpX
LIQ/WoSNmIhauBy0N1IdVfc1JdQa9GCLKPkB2ENuw7ZLq47PyPfGdVcioBInhSfdFY5lMuWJgUbN
ht93n1ZdzikPX02c70Ix9xLAhTXIFrttj19N+fw/oHM9QWtciRxlYRF3X7IWxTfKb3becRGcbPKO
kXA87ew/ZkEbb8s40gklnFOT+eFZ7A5+/SVx2uzfyL73fel9JXAxcUpUU3GZ2/CEcmJIXjA1+nsF
hMZJ1kN/JgXEq2hSHQb1/3hS8p+BwwCUARkef7qeTvs7po7nAbeaGjysmyc7wddo55iGKnYPydUy
ytcqXoFuvwcX5IRqNIIlTH9H65dgfOUlu1o5dsk+TaNzHYLJpn/CtQ1Yul6JvXaiuZZNJM7aEioK
rOFT5CaOAjIF3HwsRYgoRCio/0Ew0tr59Anp2uf8OJ9tYD8ol+RuSA4/hf7Zqre8Vs71axzT9qBx
4/KA4uU3ZnEGEDCxalMxdEit78VFUXyK5HsCXMAQ1+PP7LHqak4YiKmX7XLXG0HpUdL3w6FdBLGp
ZVZbNva0JD3qAVADA4SFUKKFC3BwMQUM67L9aEDjB/CJGBPtyS+iYqt4KlT0TYhMul9EAqeRJGDo
1na19/B1ILMngikje8ntbidUkGkXZYyhYRPcJ/Z20zbNNr4xhJarazyla74xc/0+2iNO5gTaK37T
kisTq35WrGuiSRZebTH6IkGvgAq+gEbJZabO7Qr1VyyoDP8IfNYx/6Z2tyFFUL8/15RjDgktb0XC
Gbg6r654vzATtkr1uyQ+c3OetnbgRZLsqD1xzcECgF1gn1NsNKkP5LTQvIyNeafEun4bDR899vO/
XVqegNzj1EP9S0lkIPyEH3ooR07rapC35kmbF1KpVlNC9gqmxtIj2iRDOmDQ7ZMXZRDpeqTYqW+8
Ztr6qGAwc3BJ7WnaqMBx088r9/5n6JNBXLUv50jj4XHjrG6cjooHkdGU2FBwSZXZ+r9N8y3WHoBl
o4ivk33PMklIQU8IMeQfl/gEaCUZDlbFkNJC2hYDZZaZ1FHBMBylBUPkOWDnMaZMYk3Upv9FJ9gv
uI5TMFkljLyngpPRSjvWD5fdj4xK4ieFT/doDQBGMDV2XXHLu7pTctPN0/79sN92xTdtkL1H8sYU
2Hhh4UnjwAtirSI+7LAPrYYViWh/HX26ozuVYrYadsWCZf4Bb1srTOk6sAe793MPEPhSU6at93zo
6z+lCynirpOWEUqUalCmLkHHqXTMJP1Xqb4cWtZiqymTRjD50BdLxCxNowik7w/WRyN97b6lGTv3
C/2BNqof/UIccFna1J6WlxZo7Vx+ePzxiUbIzwFzKPfTIJRl65fbuvQg19HUxUrEbps7lS0NitzV
U2Ibh1gFN6whJp3hmInXk6hEJebXgY3na8r6c8No4GjfyOGL5+08CkWoMw6C7bBD+crDFHmvmgPi
CHmL1NP1S9OhePnR6FdFzHJQazQ5H0IwCe/bjD5HuYg3ei1+yuPOJ14kZrExjEUQ+gOQndnGUiqB
bptqTnA9wl3yDR3PcOKlHYuaRDYMMPSv/3sxNzbyvztcslOAAvlAJ7vbr40wjF9opD3zs6Vm4NkF
3Wb3UvniP0ak9DTztJc6SIPV8uW/VvO4e2eY/J4vfOzMKm1AzDPFU7lr2Rl5USFosU+B/qNDJEVH
AsjK2aCo1imz6LOusjD7fXcxAdvLTrSuylUovcSTnYVP1aqXkV+jDpKKRYIKsTbpZPUK+PvFJvZL
oM0w/V11NHHgW2e8K38Gz5NZltVLdiw79lJdI5G75XU66zLbnnUkemna4xymMCzmQ/tTie0ati2u
ghN0xIKWZCNnQO7LAtN6K/FaVqHQKKIn0D3TfnlSCxolGd0Ij/bU/+qbDsedMa08NbtDrX9tLvX2
rmsT1CQTHpsfQCO9BCA/1Z6pHKNJZIRufpI0B0SebaPhRHEZSc5Vqb09WlpsGWA58KHFYCQ5p+WJ
kLY5W+eanXnrjeky1yBzJpFPR5avdTYdHIVllk2iQlloEU4NtRMVYr12XJTSfMbCS7KI4y/49TXv
fnJgxpVEsTLwNlhnW/939LS4c5TnOahz9J8tq/ZvuYjwNEThge0+7kckRz8ys5YjZA5q9wvzyNAn
BuJs3jE1dMphw/Dau4W/iNZNv5xupZhGbJEcsdhe16Z7j6TCd0KUft2ycV7jEAwQaeuU2JN9MYgq
/+CpeipxUkmo1tWdu43e7lymghduNo1E0KNFchGmYt3p+/qoCoteO8t/Cy/onuNx+JAEATX7ob0h
u1w8yzapp0hXZpOfE9J+kp7l/XGygab+3X9Lq5YiDZaNdlWb/AhEBXMQf+uvZOnSRp1w9y2eolgH
uth4QnxJZ9QF3QrhRypN5gztZ5GaUgGAy2VtvwvDWCO4v2WhW5ctzgGpJ69NFa/XZTvGnesEREDa
bzA3eWH7x4zonfMnba+AOQYOdqSa6BDBuGeZSuOlCOXwEfa9uqdpn00WxnyhO4i77bk+PY02prDh
dNfGKngTg7vq06ooVt/SJimOcFCjpLAyrdUwEgxiafveL2EQpWG8HaO2CfK1OkAhqMB57SXVx+EN
ALYXS34QApuBpFhWNHvsHzXMAdyWEPzQ7XmeOZnem1RfgoS7cftyXnDOVIZmreTlkxJlnQEQZoIT
iizJ+1uAhrylO9J01+GR1tsLhLJpe15UgylfHwohTxfhyAAfnU+nQm36Qmq+TMZ0smtZxrHYjx6E
du5qNPbUjjaDMYYLRm1TxA9WvTqd/Rn5uebuedaODixkFEoxAva0DI47SSFdjvRXEBfqQ/n3um9K
/xXjRnEP6uQsEOUO39XuDC2h9RJeIcWkrpEN9Ba5QapWJgSn/wmohuFBNVPagKkSEhLKBjPPbXXj
IuMzsad+Z1rxt2HbIHinIZzbyhORrT0nLTmeWsDDCzcdnUFWNr+PEAnCTjnAQe0nJ7pJ77dYvTs6
DOFV4ct0ST6hSeoo5a1MZxS31aew0t3vrPaQUi+zgMryh7evzfqz2ss2Lrdih9vqQ7CTVf+mdHVc
oYSjZB9TQd3hemAOBtn81suAyrnWw+tYs780ofzGbgzCqR07U0lVnmsWDMlyUHN6cyTHVigrB0UA
yIbvBIJWTpXc13mX8BfR7R59qU4EUmlaAVA3GwwDkg8ntThkE5tfaTxlbvo+Z0MClgeby+E8H7js
uU+4ImSm/dgSUirAjML+i19H+GIMyLS2/x58/lPYVz69vlcfwhVjX5D9tNdT4NbESNP9QMHRze+z
CWncfqYYoU4Z2Xb9Tb4F4cT0Ajs5QKMs74tTkd3yNuYtOUQ0R778WER1hJnUulhE7yGGaq82z212
7QlSb6lxk8UmHj7mFzitMrX4SH4i+rGt2kUoT04Hqen669nGabI+oAxjJ0GNsJg0ERhwxR9+JKVR
/R+BEjz6vbMqjbHw5YZKTUIfL9gtvENNhrlDOZSlNoQR4kdWrLWk7/d1e+USVcXQSCrZDp0O6xCU
6Zcx8ibSsq36mlvgu3HiK0hnDZdoawP1UhhwRRUYidVw/YYCPRyo//WDwMM4VyKqtORb4Ha51l/9
vSgHKXKziLZ5dQKTpWtbP5PZT+V8Zmywck6tFiarFZgeAOjEvjZGd8kAIIcJGl/Mufnhhoc8WHnQ
H0wHAiylBIs3xL3YHGKb754jOzudasCvv7nUe6r33r6PfNaVekIIuoTAfKTiKzcEfv9/Ahm9PAWr
zzNpEGsZ37f1xhZvcKzBaHAzlmVdZ/UCYNrYyOJ3gP0NAOMzN+5G85WJouwYMIXuJgjIY5HGYFCB
afV9TZRujNt1VCke6VfzeC2MXb82QWSBqpzwG16Steb6YHk+H/9j4/TnqBtyb+YxdQXzVPV2IGyZ
aSIsA4h8exrYG7Vra7Pw6HFF0gg7W7HOirAvp7kvE3FuEw5T24Kpp+P90rspQveLp7xQDgJirXbn
aK/VGRVt59r2tKm8eUYNBQ+WgqLY554/J7/l2wOsPXfVmVhVUewDOP08bTEK9J5awaoC9166/Dp0
LK/eM5+UTZT3IOQUUvbNh1kdhhTOosSs1fR0w0/KJ2gikFkDgrim4nJf64t8gTtW1Z6obAKjYPlV
KP9cT971WKYdoSbn6hrnxzQbUjPcR9IQyrkwWN/vmXhcsRUSNZwT7jIM+/gOed8ZYz3U9sOQNoJ3
EP0h1pDZ2uFJqnZ2O3Xbi1doFnxF+QWhKSi0RxYQWpSbWL++mqtALAXIp6jhD98m8j/m9hVJnEXX
6ZlHozFslolc8QFZlqVWWcub5UoZEAsYGOVa+v79so+/fhvrLmqsiH/xmvaSdYGBzeH1lE7zhrzn
h3AXQL5BN6XTWc5tehPLnpcDMp7hfVg5C6ITiADuipozAxNE53uax3rm+25Tet2139yTW6NK55FU
p24nqBbzLl6gHEUBXW54BOE/1VgVRz7nQ96hb6gzKJzpMa+HNBoJciRHJcxFfAedTL47aEEsUmRT
E3AOyKeum89Qe0Cq51mj+M4s3O7smSQx+CeaemkVNK8bGWDhnvel4sipSel4yl6RkLAhDfAx8ZvP
TbJnBxE35RHhGSLH9cOnbd0ERR5U47Pu/zG7oPtsh5Kjg+BLe2a0+TZaPh7WUuqN5A6ckoakEfZh
QPt4VZjt2x9rbc4zkAOAKZVJwpe19Yzn/vDjgw2J3aAB+U/IZNuVSve0ElwElElAUTt/fi7RUjou
5pt2jSC9S+sMzlN7mn7MLpZQLMgADd5bPYabcBdRZbxpo051VVe3D2q6SBKtwKW3QBzpVDfZjhkR
VTXRYF7djiMvVrRh6d3uUNLQnEP9hWegfxxW2vzQoDdYzHFYjeMeAMpp3xSoda4M1dLz8TcNP/G9
nMh6qkpHs6YY2fMkakuT7BpsxXYV6NEWzllSc9xdm+O6P9f5sAzejqZ1tOOWNBIM20cfx5szrgdp
iH3RQ0P4mS3mOD4KLglPGd93HHE6wLebrLmdVExdVuAHlkJGRml4ZYaKXANwfbU3LX0ktnpA/b0i
18ttb5Mu13GdbAWvHL3lusjMdLAYn1DAeM9iBbM6N3nu8YPp/aH+Gc3RvFxkNfRXLTokL34NkpyR
rpQ6THQ3TBAEr1o9xnMTQG1dp4MGr07KQubDVNgNya3cZHYGiKLJGpnNrB/gkN1kfkLatuaTX79T
oG8U/EnakqzZrpYPaPbzk/yVJxKUMZfXTNDU2qQxn8wXv2VCuxtVPADM8eVFUSpq0YvOOEkQiYNF
Y0e6sgIJeJOuhVXmn8zHuqKkKFq5/+lREV5BCCtKQY27pxeFRQbAW6lEAfPQd7pcSomwMaqxnSey
ZApABWOK47R5xZP6mImR1ctlSYcWY3m0GobD1mkGpH6B0Md84lmkE5e1qrpvRwRNKfOxS2UlvP0l
KVoXQnQe3ChJxrdsj7VGwj9+FwtpMFFdhSf6cABOaF0MRuAJrcI0te8aFiupoDZZwyzV6sszzC3V
t2Vb1Vq5N6n+RzpFH1O9kFHv6IRRhh3wvxrs446P3xbmZqNtgQxOl5M3fNcPrgB1i4DhE1tJGywx
GeiR2/5/ePlE/VW3CP/0O2NbuaTPRpO/ety2kxF1N50D3GRVY9WNKo4nDYwuJibP3e/Fb0g8AAbZ
Q1qsVuByZzQ8xg4jazDbVj2bxJkaDAWXWwoMlRrX6s0V6kLaN/dwWAFd4OFUrHNHAVm6dO/MXJCN
e8ECYHxax93/ODUuqej7XlXI9mDkvj8CJbzKr2G1oBUD/Uxi4nUbsxPe0ImTh5yAZdG73sMen9+s
JuQB1uyBTq/pmOXsVgdXY5Jw2jk/lJFQSXYBvb8PbTo4tEebJ4Kk0Lri0t8PvzVG7kDpcjL1uNrJ
LjAxkWQhnp4JtHY+VmFHGLBhESXw8nJ/7RyQkyIxH4IRHEaoA5CqI/DyqBfXkgetTRgVIv5tizgg
WgZoVcFvMGI9eqbleZDHmLCbQjQ5rBSbxvKufd7kKcpXd9c2wkrGrCRUB/YdR/x894LFyZl05rB9
rQB/CBa9mjAujPzN2oS+qmBvaoXz9XV5dURtV5NSwtyzI2tOIEtqjnYHWhZc5g6uoVoy5IGqkr/v
/PSnkza8uXWMv9jk9gEuh+7VizyhTs2afIWXtfVd4NaVOehWspXAeIxW4jPNWtDe6H023uiCQgy6
cloRfFIqyIA834kmWkdovLIT+FUD/OGnkaaN2ZzRNy9ArQiy6P3xxOkQ9+57lJCwUe2byzQrFw4b
IGv/S9QUgyWyykGxg88WcpEOttuH6Qv60lV+GI03zkfE3hGEmclBZmyB8W/N2s69VcE8hV8v6Lr3
rTqVrTQ6MtJqJUXHEJcSXvL0N3elOooHkrlraxQ0VMff9/R8MTVjT3jwRzfPLggulPwUH4N7Vtqj
gFWx16vRA13ZXFukXc60GbjTTjyxVZaHz5Lv7FLSWUf8/OB7MhBEKDvJjgfI/1tB+IzRHr1vn6Uh
uLXy5ahqGuK1FaMsNpnxx2yYKbpM+DQ2Xs3T0JSQDUPzT4I2qBwIB8/BM7ejv0q2Ej7aVZe5wDuV
XbDFGkFubePyqDOk1wDD5SHyuIZTA7iFJKt0pY0RNBonCH5YqoHefJVh5REC1zwyrteDA/0xPugn
wlxs5MlemtXTB9RF2YK9NBOe2AjEdTiSP/z7HSlQcI60qUoTpfAzeKdL7NdhLmz2w0ii4TuVWqbe
i+AasKjJx3rVftU3FdZb7cQqfS/5/KA6vR6770SiayQT2Uzyf5Hh1EJBrrJtI/7YEy0uRC55rNOa
CRRQt+6ZruTf5D/8JoA4NTNin1YzPg6D6qguNgWyGa2l4rvZtpLPZ67BiWBVWYF+TrQqe1AK2b3u
dtO67vbA/+CUv45BwABY1wc9nNJhSVDwHrmVfIYIz7N9FGkPlp0gkrnLm+k3MhlEPRc+vW4KEDfE
ppTnVoi25UCzhLvDghF/kdyD81qrgCT6mbLxbMcleM09Z9nofcN15eqDauyP1gqjwsvfGrVIESjX
vDxdCcXJu/mLSrqlhYpprxrfHELjAmzO2FdQc0cVYNDZCywX9X2xQ5GPsJpbIZZPSFUJn6nA2te5
siIoGcu1xcKSjFYE18PeuTkJka6lySAsqAn7zSk0QPdDIbv38vB8HlJAYpLmcdg6LYxrA64MMic4
kWDyC6U/QG6plitJdKOd/Ssovr36Wsp45dKpUzi0ssb5YNdUXA45YHhJMlxFPAxcxXJM6YggmLt9
qj0BpQH4wgV9U3QMYQX1XAYmX7janLWVZHjkKxw40+T3ld8/arJL1cR/jayup4m5WWJ3mzZOQLQo
ixxURU/3aMNV7ImfbjEen37h2G88ObOtjzRJxnh3aPCcjKUd5znfbFviLZBeYFCY2n/r00nQWW8k
dmfmFLPhDw9hhko0b86wh3UZ1HWs/c8lgZHLjEyH1bNtF+x62yZVLhhr6lpGlORq9Z/fSl6z3cmT
jSRzaZYj7zTla6V4YciVpTKZpHfJtpkl79RTjGtaPWZB/C4m6ZgPPwVWBZ2rVUueFrS5eQxkGP+Q
uENRFNwsl5rEMdPHTz/zwFT1E75BbH2erm4uaktpZO6spRjkzXQU6CMleleJ9MwkDiGqVv9BHIAt
6OSz/fDnQQkZesL84pz00RonL4xPcoRDwXp12kSiu/ThpNhamcb0bpiETytJXGpuRMherUezNDxR
T1t6qrFwBbTYohgs8eHSff+AaM+K0q+ciRdxk/ad0c2+bLoUUJRA/LBQgTS3wNt5oJQxfw2d+hUf
fzufJwLPVoZLN07TW5anZiHRa0/NtPz8Fy75v06wIrgF2daLv8FDV2ZVU/vC3skEfiYlXXV/a1Co
nZ7od9gyH0gysKH0nwChCIYkXln4EzYpa19O47OguZ4p0EF5upwm9vB2RLsdDlSfUqCpYBeyVzEK
ZGwdXHmiYGb3EtGbFn0hiHYnRJePlOJEojHYsJWPT49l0D/34hVp7a8iDvAhonES9G4aEJeuw0Be
kg9RyiAHuszNjQgcSS+Pxzbyyf5lNIoaZzR4OKMv/xr0by7MLAcQ4iOvvT3/Cm/Le5umkO+imwFK
SR5RuXz3sX8J992KXhAQyHn/ErEwA+jj+lf5doQ+rjor6+/OfLWGP/WKfiH3IeVkd9ayUUf4YliK
OlfMjJYQqVlQzvdRuJuA7XEhsQOc/hXeXIYNb0D+YKiJgrYHxppvSYyhPbixwNjKqP2a6JCeQoVt
+i6U5/B5BX4i+bOJJdoGuLFAnQ5tPu34db0QlkOrufSPpqMktqjXavDSM8v0IonpR6fpJHRqBO1n
vf41WLNa40HY2iaPcXwjxq3isZA2ZIiF8MRkXbcGOk3bHGg2FSnLduH640LghFDEu0Y0y132Roza
CExostSfFzQzfFqgEGb2bv8PKj6E9KxI1UtopwdVsb9vX5cX7PjwA3dVRD6osYIRYah/m2YEimcX
paiTP4TKQzcK9CZ5zOnaXN9IHo6iZJpelkCT8HUTMcV70S43QdD1aYTTtD9Q6Kg7sZxqRwSr0N3Z
ITeKYvS4bGCJLtMLF8ciVhfxQTCeUnVLVCLrAMTVhl7/O7fmMz904SjQCwo/B2l41lQqAYfqJkd7
FtwnRPpPG981iCcWyDEWl54DxqcWSGRiRx3m5oA1PjMoQkJtP+JQcYMFp9RwiLK2k7kE1djb/VQT
D1/6SPqJPvnthH98elbvbG7qBR7aJNtHciadyCmMGwdDd7l9neQKohNjVHlJh5OS/jTlo8vOtJcr
A3CLye2ttYUl1+lB0/f3aeMD9Bju599t/kCUeEH98iqdaPv+mW5ShLmQwNsQMSbmRxbWUEJMow7F
Lv14iLKqPm+4q4tjHJnW9DUMQTjWCGwBWo2wKxXjFXoTwh/U93cjGL6+BHgFPTi7XNNV/MbSpoE0
b+xnWrWqwvhZAP8q9uqoDwyhK1zNi2erAp/BS7Fc0R6hJmMZ+uwBqqE0ShWyPuD8Ij4+qUqT8xJb
eGsTkAyThUGe1sMbNdhZ6URTzYoKXISWkWyx69XCj4dXA5VMhDoaBHtEuYPg+xjydE/8zlqMeWUG
2aDaoVz8ebDGBkp0WGtpNGsKzI8xf4EFRjHq04EXb4OrCqIFXxWXvQiAHJ63v/DiXAxokmDQZj1E
csIIZ4qu8psBiGlbSzhMCxWYLEL3vmwWtzsQyBPhFCTtOh0KLNa6unHlIMpOqSCLtcxpWUbKpjWz
XosglOZltxynxMq7v0Ed1nPZaOSSQy9fWdLiQjFDlu/OPUQwduUn9K1oMWkIhgv5OlJ2KhT5u1cY
KRsDIRSPDj/kW98j/hPbkSOtyxe36aJWGT9Z/aA6Ya0AilPq04N1tN2vFi+1K551Mm4c9QwwvmnX
X1pfJ5N6hoNQQmfuulOBrpx2yYXikodU7K09CnApyTJ73+9xxMep4gIuvnPos0o5n4AZsy/Kx8e9
1IA1emGKY9PoiboLIFMRYYIoIcrmqKvFY0SqgZ7FKm/AymcaXE9pN57EbznK17iUqDwW6aBWDswa
HS5rMCguns0bNa2Soi0QkWyNBlOmF3qJTwaCWP1zcZ/0eGPG55GXePu3wlKUbPta4UelpPTLjJoO
Kd5gVyiLAFktAeN+VVAeFp54Mb0t+FJgs1veY9sHQQ/xdczYtrLNngMt9w20V8rrIIeIDVQZytWn
UmfaMxIl5EEbh74uOHWt35gi590x/lqyiLmIGxNuRYkTl/uCwHo298ksaklBCHf3cNNFG+HPhnOP
K3mVHVuzDHlFG/hSYcrP/8/hRvB+8U0igR/6pVls7av4dS3j+NSatic9r06Xc9AJR+oFXWalSTmX
mCTGAqglwiUM9bAanFSxqKEDhH2WmZx0irnSvNC7z8XZjcppMhek84rHKkVTHPV9y4XshaAdP54Y
UY7fZTOez0GTxsA74gjiBJx0juIF2oLaDRMgNV/95snPjDk5IwuTrqzP53lmNxY/RlW3fXkEfllK
l4iQALOexZpW9QZs2+TsPbRw7uWmC90DUhPDY2xDPUXTZZPFw4gWPlmc6IRKM7odeEOk4OEjTJzd
wDg+8X6Wi3pp0eMyUh1fWLrY2A3At7F9VN8/Zru5LVK2JAvHh+YvuXYZqK++nxRrlBacQqZyMtvl
5oLkc62FtT9df1NzXXyWTI95y1Hd4EZhhKjz4SJyw3rs6olmHkQJtQKRFOpDWlhuS58+DcskYM7V
2nQtgMiBzPWfY1SLxEzc5EnVL6FzG3ZLxKH5jTNotib+suvnua5wUjmy/dpP1hogwXgImCyYYmhC
0YUmOk436sEBL2kBfX4OGhXm3iaQU+2sM73SCrGAE1oDNqt4N/B9+nPuehYjy1jUUKKQ6IfYSuUV
pQ+h2fQimyAflfW3gIga/Zy3KgWXT5bljAoFH29b0ggo2CrZFP83Y4qwgLSCZc22v/E6t0JwiQmE
ZvUhDsX4rGSXkJPqQwiLcEWnQZpTsLazz3QFPVAxryaBeoafxsxFo53SyLT4rgo0vCwGHoyQRBc7
0lXSsSFUr3O9bpEhGenVtwgjXxiSWjYAxljJP5B2Y+E3e2/5WNiP5xAu68HJqhMHdJcRlxtzRvEx
NcXErw6zG98pX/JSKOa+pclr2kw5DQqqdBQvxXjlnPmMLYe2flaeNgGctigOVZVs7ahNiibyYLhq
AX95xpdsp+tzYRRfCBK3z90gIWXedXGqxBes4VnnSIYyu0NpzrKmVRbFFoiWYtJX/TzBEqD6LGSF
AQ4iZNGr3LtLE77Iy0n+iRcujRSap3u0vTG9S1DUtfbp2rY9lXfTNhe6ekOh0SCp59xtvUQ+FYYh
zgSSNlw57DICmrGdWySzx2q23gN9cEvIhoqdSx7FOmc8McxIRpYZbLx5KMFU8Jq17u/XfH9Lb241
f7Ci+qQq3wiXiIMnEpOxPNrYubk+vr3GM8hXfzgLO9vbj9UJvv/k/lXwT9jkwp0vXMy3228NLoO3
aSF66crzA01qNeC91oYHTHraM4o5K35OPisx9HdfqFLDrJhqwfeRjOXUT27835lQ1HJ+2jCeoP0a
Nw3KQ1aART1tbu7VxEoVaF/Iww65F7MAtlD7mrdj6wLOCQE4XF1BfOQq4fwsgt7KYqgax/FiCAsr
xVPWpbtM0BIWCE1/MBgJxnMW5xAMF/fAzlMGPByREeFjivblBnhWDFODsTJKb+iBHw05/ecLsAWy
7z1hDWkIwV8mx/gxHuNzvak/OqRcmTkenrxqvvXoxFK2JnhnU8WTXdqbt20Jsz7O1O0k/kZbz5jz
2mYCpSmEnwk+X64seg6og7h9tLgHIvdsATcHK7b5jZaho1i0bwnHKIjdf9hHzjsAF7imeIjVZLeE
dXzJ3vc4WPhzEcT1jzqHmyqyZQ/l0JB5lgu42RyOWb1AFSCpa5O9fKH+fDcO/NskW7FMDFu/WP2+
NpQoEhJL01b+opc5bCucShg9x467f8S7nlRCA94TsuFPZBXIRRfZdszLdfAwLN5F+zgwa/0hk9Ph
2NOIm5HxpCUE+KiQHsbrGueDcpIX2NlaPhY2Z9oZ7sLz9t5w5xgg6McguAe8Q8eGMwDwIxgFOvUm
VgoG1VOdOLQBwsn4B2v0BgPmjfPZzzB2KLgnMcnQtnIOgcv+uc0B8wYjaEwdt6p1lzU6JR8zIveT
2hZ/dD4RZdAMO++j8tncSHYuh9cs/nC4DTyPJ+g+5W0vh58/ajPmOp7p/BxCix0oUYGOpElUw5LU
Z0KW4g9oSoQa+FgPst++CvNleyDN1S1/xMiABE0l4RBbLEQMxRWYVtFnN4VxGmTXzJ/N5t78wUAR
LsETZvsM8S3Y5ijYGHFlDz6+HrApzhGMDlchbQfgX/2lgN2eww9X2k9Hc3m7pW3TaSVvX4yplwTT
45qbbOYESnyDihJqby0fPv+3G/EUL99ijL1zOcYvHolI/YhQWtXLjmgggoFi4RQL6nTTq1hTkG6H
Ahym1XHxgVyIEE9R4kX9zrt7vTyncM4GPc8Djh6xZfm//w/1eH+Jz3RHhFKjnf9XPzD8TxXrZC4W
0IJNDQZwq52MXon0BkPu7YH9p5Agt6NfoBXAYqvHH91OaKSETD0o8hIl5Ijdz+IQiqE+nFJ+EDqe
9EngnuFmcWGfge7sIfp8AB45ufMBfuAq1sCUEQfRsITg17pAe7DijDJisoHNBUqvY6L2t4otqGeA
piwPpLSvbNEUjF6tABCj1nw8t56TSdQxxXWzZ+zFctTclq9W0iZD8wXjzAWV8LTK32Dn5sqtruJC
G7TQ5Zf7QO51iQx6FeewStPVzk+tXkA1WxNc31VXyI1gCy7wK4o9XEE0tQy78vwKFwPK8mafu4Qb
y3OnX/M1BdOjqmWtZ7auW+6tWjDEF0Vp1clVyICtC3Lkweqdt9axCWm5hUpKLdYJ0feFiRPS6m7t
9w/kx7aHlnVRlYW+W99WGdWgvB773OdMrbdkXlQQwaDlBNmephRSz7oZWuWXVh8ee4MwemrmiGFm
Yds1l4dW4gI0RvT9/SJ2+irsFI4ZI6K6ej7f7JUK+OrW784RxZ9ZrG1tQbr6JDTU33IVqdf+eZ8m
vDA+CrTU/uVklC14VykR6DsNbnpNYig4IfPEhA0fttatoMlaNzrKMB8Jnvqzy1idokhEejtEp0PF
QvSQpnqB6T4Gb5TQ/Sonc7uuOsIW5JUxmzMTBiYLrcKIl0TtOd7ls0U8EqpyzHterEZK9XMguASw
/R5IDR5ferERwCCh+KTPK6zERDnheq2S4H1DgrRTvJRlO0sJ4Y+bopt0lbR8bbYPlUlZha0BaBn+
BplRkEJPYufkljnfK18dAlYbLVeOVR68iBNWKOHTjr+gbyqGsxRu0e6mvy6sLmUzk6pitAq+5NR/
9yz3ksHbPEPRVp14MEpyaLEM7xGyQo239622oCVzm4IpfucjMpQO1SfMdRpP7eFL7EJRAsanL3kR
V4itAwyWiJrtm7XCfHBze+d3Zat7KaG0i4dVEOVv2/Vxc5IJS8WdJkvXhfpYgwyTkv4Y5ZM8abe/
ukccTxCB7nMHsRDg1DoO8cF4gZ2ZGpB9lv4G3oIRxBn9WWYCWoAuwB21t58JJzA+tbB2sEYn8HMk
l2a0PWNt5xv6ACYTwhoW4d/r9428SK3jz6ylwbU7JU0KRmiKsmRvm2Vqa6sSz/JmvIcIlNcm/XiX
4KhgDOKvQ07YAoN63lu3v5B7RVsfPfnJ5QXEQlO5trQluPKjL1axfKGaUpQEHMhpt9LHBkAWMDp1
QGhdOlZxtYSBRVf7kstAjQnzMm/ynlDCy+LA/XJiTUhwayKfGc+SBlc9CBqei2R6KTxOrkDxIvrO
DpiPEeYxCGu6szbY9MfTzQzLXmJJTZ6vttS6bErSuIQ94r4rBa5osIK6fE9vB1/sCVdqbKxA8MHf
5YRZ+1+3Oav/PaJXzD44hXNYNxiUp+agjvhpsBLrWURY2l4pTnygy9p+6FwbXfJLjVPcPk8b2oD1
PUqyASDs2O/ymW3r4OYYV9ralHBMjGMAk+CueY0rUydXRdTmrGP/bP5vkdTaawglfbxubgeHNbzD
JW7YkIb941CeRumeLVnGiaIMh5oOU9tcS0nqxdppvrWjHZZhhsRpR2Kd0eh5qnNx7AE91fkZOlLx
QdIxakewOJEGVBaNSxGTpRmUJdX/neotsTpprRO2UUzaTxek8+w3UWW2gHgc4LteuTqyDq5KUpUe
zjdKLqBORSUlgv7JHT6UbOoPnineN6yOo0e8R5x32U4gNHoFf+sLNSMHVaGCpIfTzSZDRgUuYwDw
TAWBxSvpoxHgZL2HrSyYWLKltLfxWo2nP3jvzaZSay1ZfOqPHbm6a+yY3eN8tJIi/1gN70NXW8B5
kjrEb7lxxASPwFht+1T0KVIH/hRQAqAN7DDlMhtkFgThkEwPQ/9TkW/2NJniItBrpBvx/O4WvLr8
dVtG4Qh0TVLr9wqf5+H0ReYcNqP6subBHWL8EJ3BhPHuLbJvnEDuVHOlkFbOxsdfKMuCgNyvPkhe
QnsbuMndtU6DIgCl8v8JdfS5TBpNUDyc6LfFKhrg+LpfX5aJtp/esxWyXCwP6/N+pTT58otkf7V3
fiMwLxOrEd3zOkkJ+HfcoKVePK1H12XnLI8CpIKAtj5cV8HRxIO4KAGDfS6L2WBKvJNXYLY0SSj0
geralhE9HbjIPBZ8qbWBUAlQSmY91y0iHlgnA0NKhDmcRKGUhyXAajhqC9xyQNEsQnysDSJSQ0/3
x24DkmQny8bo0qrYh/2l699XUR9GjVSdUqYpy1FkIoeXzmMLNe1nl3CBY4wDE/L5VEsfWIfR4oxv
qDxpNZ4gLRW2gmXPHbeXtxerxYLduO4n6uw9VA6uxR9HH6k8mZ8xKIArJN5qaLcbqhMrjxSxO22D
ANx64Wi041IdnGYkNNZ5ZEMmnCvgTCLfXdjvV6dvUA3sFFbH5j0mUuhUfjQz0oKv3Bqlp2tND+ps
jzrYXfz1FnpyiTg4jtieM7JazasCCnzxbz15bTKm8Ed0gE3XCBIGVFamF96cMAf3yvFJdzsLw8Mm
o9gsMfdHcwEWZjT2f/OnxaOY1YeztJ7YZqqGEPRU0W12GJysiHyBSQZpcOsP2C7m9CMVyLXdruDP
MSYyAbIG/hu7ytPBD5OfnhUkEtHovHLm1ym81e/QbGI5dAj/1lllliEqSu9bsbV+ibNWthHIs74y
ceLTEc3xez4mSOCXfhZNsNnd2KsLaHoQHgTHixfw1/oJxGVkr7aEWolHiLbQ08Zyjj5fZHAhqwhI
tkvzYYpRmkoWpvAIrd5DDfK536lhCAa6T0AYQ6hy3ETiVaEDTKYPSuqvU6RMYwsMqBtV/Yg9gv6q
kGRZJTb6AKFe8si40+La0Hj6rUbsvNq4DgMJOtjSKKd1fonfw2BpOwP4szXieJMU2ZB1qS0s/Gun
nExuj0ABQNKh/jq/uIRegkaIc0hTbQ0WfhQatD+lXQ93wRMLVv7gQ4DF2V7vPZlEJYWhS7I/4Bxs
nhoPk+u7Fftmhv+sqxH8mO4bM8NIh8CsSDa7EBLbMlGxj4FrnzIGvNPU31JL+5h0D4hIdj6trCTu
4L1iS5cW+qSlpsfDfZGrepdoGv+V7GfEr+onTdLVDuGgJwJzGHFtnU5JUwlYgFa1y7ek3z5rMIP0
UHKw9ucdpqdx9afX9SVWwjzCnvG2CKb1i6S/XCvmazTAbU5P9B7gqiPV4hIZYm1mAHkVw5Exsk0f
F/Npaa8ZfJ99r4eykZfxIcYPcug2MkIo/3CQ2p9d+GbIBReC8XOS0OVaySWmmSA/4zRKzUQ7oYSv
mTJkYCkFdDgFfCR4o328dFOvKghpaC3ED1G5ODLPtCtgjjD2nc1zGmastE9BT8SGx8M29el1SyB3
htC3yBpsxx5cyaWE4gnctvHm0cp0lpZVQoH0/5Fj1J44r0/UjqwXWIzgNYgy7nixygslXvhhk/55
W8kej8qsD1dbcjrMRfQD3zaUEL8dShH3CWs6y5QQZ7ffGs8JUIMlUemnVrokrUoe9scoDrGIP9Ik
7hYYSIy1cz01byi6h/25tJw2aM8zrIiFRWZ4QSKOCx58wVU4XJAyT/vKnW5khnCIRlALsbKmura7
rNBpMMvp/G06/a71ml98VOT8jPD6KTfoQgMeHezjLvxQVsmoeew1YcwbfFUViY158KwBw5alcM7M
xSm7dSLotWv3U7nfwBIx22vrv4PEl2HRSyrJRI/7Y7ofq7EN+paY51onCiU6ezHOil/hG+VzgNnp
gjYfPeyViDykoHrwiWvk6/gdvSr2PPT/giK41P+NAj1Sip9/VvJJ5an89is12iPtiUGRknIcDDrZ
D5cgEKPybOqKx0AESesJXBgNUYqtB5sMhzlozu4+TvBzDtoAlFlFsDLOY8lMupY17GkLD9a2QLmf
3OzZat96+aceHcZu46OyfNu/N3+7rTMlITQecOo+RklqzL2yBRpkn7K6i0I1D/13X7bHa9vapYnI
wCmPaRFKD2kV5qKJWTvIgpVkiylAlNHzKDWfWmKOmLcGuSYtwz4spXRC73JOcles1OsXrA+vwTEO
LDiCHIR0KXSGuLdQKUjtATj4NGHu536kpsVSqofPDd96Klf7P0LjpHZCieilCPWtX8ZSXYjHiwFc
UCIU/FQYUSbWtLBPsapZgHL2OaaEuIhFWtHW5GxzQ68D+Bh7fOUZZXKsVOzyDItvqUK0sAJCSUA1
/csy7rqamt+2zXWl/6ybaN+WeoXgcbejYpFrcrftqaaA78Za2oHftZMtsmzuqrsQ5xlc0+qRS4kf
XhowFlJ1FCKfKARs4RYbUZTs+d6+Gn87sCus5Wg3pCYCom9MHo3O3ukAlFbYaoZRYTg84h6QITod
OlzSdX0UQqkwuO+ZPMT6Kz2tIJ0AO//qgDRkgm1OXiRpO31/aSBELM6VCfxZ9Q9RFEp/hUxVXz86
NajwBTfyYtVMdU8CpLTgc6X8n+pEFkgMAgsRsXBLIF6UQYiwTXGLnlVnUYHxTr9ZTkHyc3srfuDX
pzReE9eqUcyJohmYC+0Fu8ngYeVTW1jpC6K1aJJDyZFAV/zwmkl+UWhbUvBd5+0tMWNo7YtbefBj
nW5VIH1Y9yPGnnGAxxxvf30tzc+AvjFSPiOG8MFV9ewHywut+NZuslJKLpXImENbaWd1lNj7nTZD
nY0KPHPhgHG0RnVtp0Tf2QB97ryccUEAzROzPyRGhzmEzrOFk/Sc+U4VlY+kKdlKCISvkBwV9i4M
YZY4Zeo9AXjINssurnGpQlkfbanEzgZ/q9xmC8+B2JWd/xf8CfJTGTfgRHbrwxhS/8FmHGKqlvhC
dz5Cei6Vexj4ySkboW+BkQ1l+oPIpgOBkcVvNX5XROuycFBNiXwoB0wjsXmZW9kJR06e/tysFObn
+Jivj8judXZbi05hkre3wauYIrEfU390QcMOjCl7BQHDbSshua5qMIYHZj+WDJx4m5nzLf+INzI9
Kg2g93K8WiBw/Fo32fEAYgch4gQfzNdHlMwqG2Zq6QY6CXhw6tPEkKFoMXELTJgdExiuCKTe0J0K
0oaCnaTbVyJ7UbGr5s9Gme3iPKAOUY5eeYtEU+KR0M/Yli8bQc4wRU90MC8k1bHh9GZNXf52gJf6
mv9IdPYywJvVNqWUNknPoxgo0ASIJc/+3XwKVt9+Lt+5BiGaT27HVbIprFiFHoPNyhn/ty3Ize9c
20ulJP6o4ErafDHaceO4pfNx2XaPc6+yl8x0m9GFKZpBkQj4xYXWxrPXXkpwlM72cnPqi+gb5AJ2
uJqlrMb6tNBypXEA6jselU+pfz1tbUKNT9+B3jO1KF60jTB527eQQE1de/rM2DW8apX7y1iEpIcg
sXGPo66Oj951uFbGRYfniN+9a0zQRwr94aLi/2+WXbzAed416Qi38I4/Ar+VvUOOxgpk2rW082i6
MWGKRIupSb+Jol0SLHf5kePezK47NO2Rs3uhrd7l/55gwU+OurHXBT1XxnfXPCu1oYCBgB0QdjHr
qmTTgVNLxqs3Opk1L67ABUHpdIHbofZAfNqYpUsU0vj+6jmHyHjmdPx1kmg1oyEZ+sncj6rYcEP9
X5WnmNgVESxgpalMOLTreJca1rCTsjQsnEtRp3IhNlek3DSZ8eJVYCYuMlL+EuMokitVk4sOnGIW
fELqu5Nlrdt7aI3s8X1uT2418oTpR2gIJL++F4t0mx4eFL2EaBfo4FZRGNv6y3PfA/T2HMBC1Qez
PQvKQmwsDBR/9zu2/Us0pMywTqx3jLGky/B5h68Eaul6+OCvkGD/EmhdhF1ko4UHUKoWNun/I4e1
44MAVctMk0Cw6p0BGFCSaEja3criaKYFYDDaLxmsBGomXNWsL8hWlcHIIyqxpxE4R3s/uqom7Fmm
yZHqHPZuuVr3Sq71nxIhrRMKBMv+6RRcAo5TooAc3sgInJvy/a165gOFQ40EQqZCENpzcQ9U6TZy
qO/Lxs/e2mLzIRI95I0qVxMoqmt2mlb4i6L34yAc2hVyRGCYPnbpQKtSzyS0O2CwIzaap7CvHuyd
4BkhTFyP0NlD1wDnIH4zROQSQzzIhhmxjErNctxD/8m/tDew2XhS/WQoDNKXqMXX+CQtyVZ0u6f9
ATTPoicBwz3SPVPhMyFKpP/NHjr1ZNzb2re+7E60Xu+m+w4SkPm53PUn7k4YvAfj+xd6NN573DXa
KKtRYC+htst/vbb/VvqL7qqvtg6ziWaiIRvzSevGSCJ4GVhIHkOeGF+lO2CX1r+ef6Q+7r0pBu5c
JByXjl2K/ORGYkPhRS2qtoWHv2wee0/XBF3rxEmq8BoVm/RoaBzuxUus2DsYeRcGK1UOqvUYMw2P
SZ2tBv7mYqb1sUAblWxZS9T3qpH5bnmup82f87EC78lfh3TeRlyaPzZSZtVb2aOoiNBbkW7NmReQ
szEXbESFfWfFBYNUApR1qAxIvnZBMPWbeS0GQqiQ0fWAYaEZtZc24Ib7wGlw/L9GUbO4gT6wK/3e
djVeQ2w5dCiDLUcSahUknvZo6OmVQ1dglq0wPcThE7UVpfVhEj1Sw/GZHNqoTvW1hO/ZFvII+ITw
DbAbS91xK9dmTTRIbzX+uaKzILkPXnTGHwAzSV5pAwtqa63dlg7YTy5cOR6zAON52ntjp4ATUCgR
/KgYnLcnpaTaayUK/tWe2RZ/6cVvpIuMdCQ+f9Zp3GB+mbanbSfVwWTtC15BmB2XWCEoj/rDudEQ
J/iyAHbmfvGdI00ppOCSArvDWiDAC2yuyeyUgG8HlKobq5fSMcwt3bkWq5FsDqUtJAbHB3nKfOtG
bLfxX6FzHzQgNRFIH9FJp2me4SH5oFDNG+YeZ3dqtuZq1aab4GoTL8llSsTTAD0oPUBqJFF31Gbn
xHO+ABUA88tDszMWEA/VuiAtRvXf4kJV1MX+JBR+BylKGn9ZKaxv+lIMkdx3K7VL3td+NXUgRl/l
W7oe0CMJLErtnisT0icaqq4Dv6+I7nxLfc1iu4YrwrItbcnWGJAJENYEO7PaIh5IAtU89VAHo82o
X5zX4yptS3150QqM51Cf5iAp22KDYRY4tqLOsXUyjY/jJ9SCLBBBrHZpOGcJ5bg55Un3GVmenNMJ
Qh5ffE+6ZJNjxrzklYHlrr+tmFK1fpKl/g9sneva78UxMmB/fMdPw8lxQ50+sv3il7ChBTRGI8G0
RXiovMgS00rf/zQ4F0aIA1/5qkaOkaOl8OirT9hMIKaQPJx7whusxxzLxnTzBE99MJw6KgWvktLp
iXVkPUpW0CSYYm8lMmkTb9TpMALve4cvJhlcLhlbP0Llz7Sw2aMuoL0Tq57rg6MDAxzN4ZU49nLA
xQNVyOJ/bgV2Xv/a8nx0tEg48iysNRMA3E0TCzSY6CoSSKxSFu018CYKH9PHbv0YZzmfegdwaRQ9
zR0yo9bprJoxNIPG4tIflTqsni+Ff1gF2uSWFaxyv3M5UpcnC3gh26gQ2rnQi5QlXvgrUDryqTVu
h/kXoUH7Z4sNG3/Y/sH7uelx9nsoZtjArD+HKYVUcmOw86DtdjsYmUIlcEkrSe2ezOFgLKXOwA5M
4q3/7OAGG+nk2IwfdPPydNv4BMD84CdtQjdN0rI2dU46AdkB3u61mrzXMJa4kz1jmRqWAJ4MDmtH
4qWJjoM59dNYWY8UoTTsONB4ErhLsnV4aCNtSrfXXdvbHXKAgGZX22MK8X/hIUThOdA6EKTObVhM
OTz/SGdlcY5548zb3usAR+8gMFrW3+jLXntb/Tmmm0ely/aNi6MM2d1erEB/BBDo/mYst0wHiyxg
Q970wgbgZvd9D34cVOWms2VC/jc5ITHWIx8cRfcVCuKsT4KSwrh7NiBozA9Mx9st+FrxxIiphS1w
JqE2GqvrJ+OsC+8C+lTqaLsEfeP0/VFtT/BuRxGFddTSzBByw1SB+rqsCWmzvqXI1Ah2LI/ZTai9
6CSnP172UmSs2JPUkVPyU6QOtGZoFLOW46Xkhw1+my+04GlZ7tt/mnrl9TsKmjcgxpAWIe8dhcbr
uQPOqfjO3XC2i3V7cFkABipX8aTQ5WTqFGM0Gv/2gRamCgnNKK19wc5Zj+E5mF8dfPg938jMUo/Y
5L5NVFZaSUG5h8A0IuTJyoPzKIYqlQ88sm5nbcMmScpmzk9zgs8ZtE7xCQSUyXWm0ebQW14Eryfm
Hp978iv0BrfR84z7LgHReQAhbq4p4CCBMFoiBhbQvPKXH17gYkUUHfiTxW2XuKJOCT6qR385vbe1
p8wdYoySr0m82hCn4V5+WzXmloXi2ZcgLSV2OPfP5M903DK3JODeAGXTre7eXYJsh69u71on9N1A
gIEaG6d1SNW/HQRVoB4IlXbUcDm9h2HDR/xujWOVfiKaEIHtO1MxDIO/qqRBF1h3B523XHUS8aib
zMWnjKA1+pA2/UftLN2qY5YR2LrWPCrwigfkB03ZFB7nUgBfYgqd4BsKBDabqjf6CO5pcklmeHhk
QXSaFiLmL47u+NcmS5/nRXpHznXlkTqALc7nuMKPqQpGzuJw4D8QxDl9oCjn2u4eKAtOxeEmKgQx
uZKGVNvulRLT7bqgRYMrPi/Zvt6FDVrihXXDvc6HY7b8PpoOwhT63VnEve67ggbAl+PLvjwWo0h+
3gYpp4zcMM9kW9qnx1MI8PHr7w4o0FhGro0BVkyVui+pHPET87zImDo6I3A7xZghoAAVSQ7IUh1I
bFaPMM/t0tCo2gJuzPgVZrw3BbbyKZfPyh244S1BIoQDOPebUYgsAvO/h5Xn6g3Ra70KuhgtUIcH
QMyN1Yh6P4SqqAD1VfrGiEMWZjKQitmwv04i8EVlEJjMVD+9eyyX2GesK5AVUr038Z+3vTzqSqEM
0widk9hoA0fSkPSV5slMhUEv8rV+F3OOIQFo3QHjbILV9EY/oHWJRADAZotw7UQy7jq09dDQ02et
4jiedKzUnnWk+Q19R7S2LjiRdJJCIY2TIiAQq1jZcxkUtx/OVyYPpqo414BLZfsgvCbbRwfHIeRj
AV2CCKyFK50lVtDXLlH5UaGcOhkyB3wNhT66a0TUVZA/sWABnK+A84+aiS4pL5ujQinX2S38hqc3
heYIO8DQVNwralNwCIUN73FKZIdeoahueKyop8JLn6i9q1XMz4yC5t+ZsPRXCNqlDL86m5FskShh
6S64ysLb1Q4j8XjrYp31OJ3Tp6HRT/HHTdx61a5pSHATLBt3En2lz2yzHq40sgbyY4GPt5mtd14B
lZQrPnZGUE9LiHZVsZJoGQL6YqovNImjwFawbRAkmHEir2Uk0Icgdc+Bw/LSuQMAWdMkVaROCcgg
ysb3Zg0kAQR5qtxky1cZ0+FiCYycYgHRL4gTrVjrpEJTSxILlzuZrufV3+eDnHPTlJSuXyE9qdBO
//hIqA/ZNrq2EMeqSqFWuvvKatO8P9REU2uBd8N8e/5ReS9x/3SVpEwKPSvdQDKJmaIMGvQ1rkQI
krlr4DEmRdC9jb9aX85BLRntpogOgAB3T4c97qvLRD2A/MKcI6iINi0WOg9w3JcOsKcFHYDqBa6R
BkDS4w5FqdThXOhE/sY7omvKjl+RN3XnrYbdvh9gMY4CFipR9/iegJpipyIwF86VURd0EeUxpqHP
gZ3/7jxEXCcYTIzpwdsP0AkHsVPCiGdbX8sOrbgo96zmL3CreLrWA2yNua3PPmTz1joszev0xR4U
DErlcMlXthX/7HzS1xKTVoQuWT47arbBVYeDEFbaTok3MrcbZ2KPcH7mhNXsTR8xU2aDxPANuFEf
Awu3kJyRripeCeQtHnubrKFR1PsE+YwNjE4cPr7yHX8aImEbCKV5lStN2hMgdoKFv3PfQvcfBsrv
0fjdjbU6o6xmmXZLuz3qFlKEaJlF88ha50ULI1ETmfMp9LAZFPlDkfF3vr14GWM0BR/jBaC//ThP
yxMEz0LABzJD/Qyevj+ogU9MvRsf3O/Nc/g/n6+MXyhxN8DGrVexpuLowS6015BCIzUC2uIWkBNj
GdDlyoZH5b4Q/k0chizygSxN2prtfS3NUCyOyNNwSxQc/QQc5uXLK+vcx8zVyJSQ+0WeNvdv2ekD
IbbPTLakEZc3ZujqmhEScaHyAC/ID0fq9BjcuvVvn/5Ky9y/O7U6JEpPCujoTF5WHm5P7ouYkE/T
FmMnRyUdPEeBaV8AFQVfZm6Say7jijhsbTuhUB4vYBayN7Tys6kNyF3rBvx4EIHJB7UKq34eOk79
HKBWeP82W16r12inAQzdltZiWgDGrrD6mfv5/YUjJnEDm+1+e4TIYFjQp6+xGrS/sWLK/1bdQLaX
YOs7LSud6uEYpQrkHunM6IITQdbpNxTIiUeMOvG9b2dfJPhuj+jKTIHWRU7zNxVEx94IAa1wc0Pf
HmqgxkobsOAaP+zCIU6YtOvue9y9bW3y7bM21Zrgg1AQGumBHjkb00T7VuX09mHsRVxGZTTR6/ej
eFOoHjLlilf82HID+4Dxmhz/MUm8UgbIJO0cAyvo9dFypjfZX5DeRLvwEGyGmYaTTRIgqLHd7uA7
Gt9B3cFajj2Wj9DvAfOLYMWwdULAxlcuYM0zgO4Zg+/w7PK2EqchZKd0RBBdHBodon9nnxRNduNS
SgZBERftUUq67xhpALvNmIHHxEtQEhwwkwzrwmm2+Kum9Mtw96K5/bu4SwQ0iiQzAYv7eaG/1vzX
UH/Sub7PTrgbmGyXmkQie3pzArKP9y6pXWliKp3jlzAT1uabMipc/siEgE8swxr7AE1tbc6QEm9E
Z4RAPjsEa68GMXcEADQ3zCuYzKEdJxb2dgeenYg+rqC1scdruEycBpl88UJNpviLUcjzHBeK6M2C
BwLhGezwfJCU9IOGEry49ZcKI3OOFgn+1sj3X0LZQ6pPfmWxFV6nLc2FXesf5nTtrj0TZRcYJASL
7sYWKCM7mD812RLLSW8DLoRDV4G5yW5/pyT71NiQNk3jQshyN+rgV5CaLDoozijg2I0N1WN60V4k
YFNiHXZflXdbBA4fC6ImC0smMlDevuL7Qa/zbJt1hJH1j1mk3ntpCb2YMj8yRy9TBlWNNbGwj+h2
HbQWHRuIg1ibo5yNwg9dhIv9RQyDaf8lJAaumrM/nGeVjjX4jgdus6DhFtXTTS/MaNv0iI1n8cHY
+N9buQYWTDhPW/mb0ThAgWpNG0TZ2JVEoFLLj5YXab7Wi0pWHuNWw3Vj+viK4YeMdTLoHkTthNyx
LxJKRVoqStpfeIqBo3q15h7KqfGgPZhXkLQYjo/jVM9DgbI1oX3h3foXDMSpVgZ5ZJlJTFHlyfoL
um3uFDyEddvlDx6SKdp4cdrytvykNPE7qdq2huRmtm/klA7oHjWP0RAO5dpHtxErb58AOzj1fdvS
TQisI8y2bWASUsc8Mq04uVh9eikUY9DgFeA/lwqTXnmMANOOhocwhuklcKqzaroNLNIurGGNsX76
PGFLOn2tA77GWL5x/wft/yBTJY4k9d02d+12bMgfLXFEC/DWpvXvMBzhSRC7CyJ7DcNEz2yb57kT
91CIlWJWwxuS97q7PbSZmeRBN0Kv7PN1oueetR9ZCU2JYXYkgVvPYnAADYgZi0nGcGOtKBxxFfCD
FSwQYFp4y1ImS3CakVcdB1TRiVF2l6CwRrJhpH5xB1dH0qi7dIxV17mmMgzGZZm01VBURfURuLR+
rfWQRrfYVBoBVisfNrhFDaFjcNGHCEt+dFAcG07wQkU+IEH6P3captP6HgDlPWypnlKlKtnItwvL
YGdLvpEdaA+mbscn5mLknsQww6QLukPbTDbF4k767CxDxBbi1OwFaUTQdVFOslukdusZEjR6FGe/
zZP9EcStY9DRYwieutkvhEK4noAsMC0V7/X7b8Z7iakBYH62kT4CpOkfNwPtaQtf4sInzmjLRIXu
Yu/14aZic962dGw7QiEYpAQ8U2wefGHmAUMgVwhOQ2K9NCH2tUUSjtaYuT9N1OCrabMgpKjKwLE6
44PgMQ1MkF3mVPPWtkA9CjIDhchcDdxbEiuIiOqrpZHGr4WCDUQevsCNgYu46lTFWnlVOu/cuJgc
Pv5qZGoKfG1QhQIrom0ddIdYqJBla4LK6v65Of27VUt09QVDUsXwFY8z39G/2PphTN2z3jyDLdT0
uQsbuw09M77NlGi5ZPmfDBCyNucgnT5JeJLWDJWbTKrLIN+Ua/grE5e+lmpZBf0OYpTb4Ehx5P9v
mYzKSqzbqwaTFyuy01xuRbD6wqRdqQj55oz6i/sN+7DVdjxGy9L7bZYJyRzDq8PJe0GGLTJnglWJ
SbV2NSvBtzJys6GM94mcb4MwCZdWG4G8pC6IJcYAznmkoYTQBBVI9k3Mjl+mcrpeIY/JEFh6gBCn
YAoVbKnNLB1eQmjXLMJkTkiZk5qgUNrhija89QlEwWrhwXQWQPgr7RpKg63PQ1Fn88KJj3wqXKhE
BCUHTj/yrkytDC/0CR281DLsWboAVDkMEfnu5YI31e9CyVczH5ScCAW3OqPsUo77Ry5dA8HbT1IU
cU6fOsAJDHMJ6k55J9GEe5nzyvuAp9JXY2nE5DBClFkXhvv6MppBiGL5H53BWkBEDJwar57+6jBL
fmegUCpi9Vut4Hdmml6KfVO9WolkZukZdYvFBFTglm0QJXWudLjB7M6zl6w3vOGuo51q/8pb3CLJ
+RheYo2NFAXNNRIeiXisJErrSE038QleGKtdH0OY/PxozZSybCgx+YIrJAZn8s2zOD7y5MOFIose
Bq6Oe1qQTBXks2TbC1cLalg+Ja8D8NGZUItL3FM2uA9a7l4iOGV2gvL8VrA8mJwfVv3p44RYmM17
1nIy9LmzvSsVK7FFhjjwVzXNHt/MoUn/W/PxuzBYPrUZXy1CjatjbtUuM3sMAdi0J+lZRA8X+qmS
iBv7S1oCLTpg5kxdzB7E6xvSlqcUseJM74PnpUW9OXKjHp49ZSXOLbK6vxP6Y0/XrMXq6U3n9FpO
N7+9JB9QjD0UbLYP3SktX8rCC7hOK2F8cj1r7DTXzuUVVyhenROLK8uNfsIXYfp7aTa4DjqvVVqf
1sV/WmFOnHoyV9ABZ+HvToGVPPeBT4MrPERCcBq+sdt1jXvNCDlrGTclahTgPPa84Gvf0ozi5diw
tD1FeNvZ9XUtqxBiGnB1jlfc9TiQuijiGlIqIPK9mK96o/jvOviaVVXRxFjExQsy6Ke6LIQ6WbM+
cxmMl68dix2T1q5mtrwwfBdxpz85JInvJfXnHuH3ILtLwvBcHWcc+YCpu3OJq//Y+gnFbc/jTTZY
bDADS92XOGtaWEh0rUbUjKGMO55Eqz1552n99/oHYcxdU+K+YdMzERF1tUXkP9jwBp98PHdAmYw1
LuG478MQSBDOImcUti+hJhv/UkX9LRRWT3bjxYy9F81Y/87nFel1EFUB8RgaOj6fgTUyLRAOsk6u
kQXBMp1QxfSsaAYx/g3cvfvNODHRdKtIM0r6+9FtIzET7eea2WR8/+I7xXsjta+gfYVuqD3rTNCC
/zcE3MInXyMfxVzrnZldNSur87JCPJwKW2LRY7eZu+npUyXWg+0txO/W7P49S58eoltWCJM/vvtU
fj9Z2fOECkXtc56L4AZPZGDNN41NaD1DbKIaIfqQ3YbyWtGDmtjNGYeSxCF16sGhmktL051/sLyx
FjHYzxposw2zkkw5FlS+5MT4MhXhEnS26kJB4VrfhP9qey/LQfnpT6YXu1TmAoVmTuDx1eL3K4Le
lxVvBfni3oYdPKFPWL8RVKREaAKi5TpxZNbuW/LZpoG+yQhe25QMYv6waK5SBgOyNLM74sk6kFqj
11OEmgebTvBvrZE086HdiJE2/fVCyKRij4Bvl3UHY6mQ7caPhlm1GCiuuQ4KZvk8ciVKfjl6PBvw
13z2+4ts3snbGU3p5D+rFipu4LsknVzDa9l+l78KQU4ukrwpVOiSRFCp4diJVe1XNmOGJS6puSXH
1ue0FZT7BSxEqAW/mG7+bfPQQS5oKXJSDt/Jy8xuLyQIFryv0IG15LIWUyHIWZpW4dXkLo6E5pRO
MLRBDfWy+O3CbKxKx7X0W4Jm7oD9wgWVOxcr8notx3GFtvOrZtvqIgsb+L1E9FsZXBgnqQ+bXqX9
rYWbmypjwby8KMxgqiahGnf6y97e1P8YzZezc/ltFG/M3iVJU6dQsPZBpjQJVCuQ9QDWrfVWcQMb
GXWAmUAfP9kQvzck4Bhdsq+PQeZD+vxhkIDKDT9zDRoUeWnAqN1zN1dFHTSSWbB00Ho3/9PRVn7V
0JMMDNMcHi7LShNSCaI+JXnFYE+eWAuSn1NDGryEgqkd7FdEYrOdTiwEOYeFww6nAYv0WEkMeOgx
Nw2SFHWYWj03K7i05agScs2CKUkmHIxxRK350YYoxhe8utwaRKrqaoY54e7OJcv3Yav8OP5BQqTh
Xwv+zOtunsTlPpzxBtcI0KaO1TG53ZfO2goGNKWkk7a01rDCueZ+EEx60Cf2jK/Xdcfewfz2Ldvf
QnlVGc+S4j5hm1GxbfO+PF1R1rLK6+M5cu1HwUXh550Fv/whKbDpCXAoHS6B9WyaKOyGJUGtRA0J
ggGq4RNY30iArVuPJrcQ6Av2UbV1f2PXS+uOIv6zFfoBFIqop5nq1/+jNmbz/lgQOPMOJ7JfKRHD
KxV1jPiOoTsYMADQDlwvhijIcyGu/AtP7PGGoezOdu0nvYtT1Pu9RfA+xxxdOWLsBWsodqOFfo4T
vZhbJrTMAt/QVhW/Sk2CBuR34lYhjBA1u3UUjkoDM3THxzh0AzNyJHihEHnoA1F4ZhnY2vLF9tq7
0fnFup3ClWVOozF6hTiTwjIFOjV78LgsRIfdDN+AwwgZzeWytNMAdESJm0OvguogEojpFCV9Eoat
OXVhS15HPv3Np/sx84KT095CcjkwG0Vhid9NbXcfjYKOSXjh1zupMz+6ok7h8L3UpkZAc5a7qRrO
8agagv9E67J6LCy+xZHunOQ7ib18rAtTYPSr0ncC+CTqDxSEC0vLCmfJe1OCIlbQ3WEOoSINT7zf
Ci/cS+Ccp1NntqJAqraWUsqD6mg484hu0rQYkq8PeQ1FNMeUTSisOPcpPGWfEsRho44rHPYZPauI
Aih8oE/tDA3uJOHREDY0VOTsLQHNEknXIdI4wM+qKaIJLk2ZLiBBVfIdb0tsFPn5mMb130Hx3WZW
krjYbe4vVfnRIWwhVxoJUBshSLISNSGODST2Thw16LSLVvK24WPncVGytrfcOK7YRMH3TJOlT6tk
fya9uIgt0nlaIhLvN4xk3QV9oR+scMZ5g7tbDo8mhJTGJiQHod8G37NPY+wQN0TdcIiYmTs2o9hP
qTzbL/8VSy28YsrrBHdkuWt5ZwErkyWil82h9Z15wbK2O/4ea8d3JQ7VhLJwfd52UArftbZSOlDt
gv1xrPmTaGkb0ZHYsHKlBwsDlNEDblwA1zJtAzeJ8LHCWh6mdYVbbxz7F2XhKAxrkqGCpKCEEKgB
w5NQd3KfgaeXuyeINI6JDaoetHHlHrulGRCGI9qdOBmLAlOdpXYeWw2dG9Mex/vCeXyjuKv6YUHW
7kuIgeaqzz6J4aDSlNdeBHcDA2+jMyRYNCLw2Q/PPHnlvnmmi82IyMlxAwXhOZZQzhBdLqoGWc5r
EkhNb5L5CfFDYA5Sa9zzsH9KRNb8p7qcnzJWguHcbbFHXRrLecFvA46eEEVOcTMNQ4Xu9htd1Rps
wpXxR6PaMh1sCh9G8NPpDDg/aLT2Xhkx4vFzBiKYIsfhzZ9VQ4oqHx5vgHw2/fK5In2Qxd8KC6sm
6F3emh1Ywk7SkLuc13+m9okIztCKzNewmeLnC2C4VlIyBikp+b8LI3HLlHs1XOkdU0VzK8iUjaLm
/mwfxyN3tCcJUfAdnTgGFCIvzUl9tZJbXaTiB/g7eQeKncGrwXkT5+9z/Ik1EsxO9Dc2TPTxUqXD
G1lozM9k64EWpUhN7qsl84ErRGFZ6Xg04PQ+9BGDOZrQnxOOAiBFqnpcOseZixA02x5Optgq21xG
hMMPg9yI9xg07iPPKYSALSZyueO8Su6/2XcFfPHaZXFr08RFkMkuNpFsMG3FLrf3ChRuktaUu+QT
3K3l4hvr5yFZ+jAcduyCm7n5IUPVGnSTcQRIuhQZM1Lj208LzkSywqc6ZnAFhkPBUVqLItWD4X1J
1OvNe0xgTFF8PM6DVwgCEEM1Y4plYnGF5rUmrY92s0Ocj/N9FOkKFgqQbDV0/6CY6td7cHGu30lx
pnTvZZyCdNQ/HMzB+Y1qhMQxDrdmViMvslIq+cm0vj2jq3YjjxELlFx12frygIbijIj1RgAO3stP
YLsGbVQHtHP9F5D4nMgJ1KF/BN2PQ6VmFpLUjjQNfJkihONC3SSOLlwVDFHiKcFZY500dDSqvASC
utHDrDOjz15VwYtMkH1Sa6G2Y3UM3BFEIcdvKFzUgipWWf6v+/RbU+hDcm2VfxjC0lc+o7fC4+iw
foKE/hDJYcqZkaTNHwFGFUuQehs9iqEj3ezthpFBnvNszGxOiLh+DexLZoK71DQx32S2k3j9aTfs
mXRgfY6PcLp5VUklQ+dSkHfY4I4CujpsjmL2tS8ksXsG6VnRPZcHolIDnKEe+NO6MHBdV7+dWo6y
s3dnzzXMuu8UHZdakkRi6xwZaP77TmQKREbDw+BfnMJUbto08mp3n+B8U5EvgarCfapj5xB2cmKF
iKnUGnep3Iwnl6qa/BsqKxxYCGGMnJJnCRU/OvixWRT9wlCW9sCBLak6R7ALBW5Y6zKif0dRKIhQ
nKTWsFtvPNXXkC+BDdcrKCs+iwj1QYFXg6Kr2YFfamj9xo3lZuB8MzcrUsCWLq1/YzdkV0LLC+vm
RPhpa8E6prgcH4d6+elAeRNWwuNmK4CxGVD7DfaI+AOXoJ28X16INsXKn1VB21q6wxMHj5803Vqb
SwBS9rjz08dtUIlRVd7LGdeQR/AGiEb6RX5LEpnyHqU5j3OwQgqX0A6A6Du8JPZ/6Ih3znSebiXj
rZHNIW2PhB19kIkIZeafhERGtVnaCmSPmKFFDcJk1UzseT5OtVXX+bEdwR7TG2pneTxVTq8N/HIp
AzlQJJf0thP20fof2Cm0Rt+TFK8jTmscafNQ+yKq2BhWKFpgk9vMHTOVlsJ5CiaTKZlSH0RRBKGX
uOHyt5JZl0kIPy7YrdK7Su1GpUM9dpewVfquAg9HoY2mgW2fwT188O6ET1glKbvn4hJ+ZCp/0Myx
fMz+HbIdc2/bvyB0g0OjC5V9CSiMV43XWjhR5QhzMaIvVBJgRwkwLeK4wUtrcEYn0luB2Rz5OSwv
ayIweN+U4RCqrOzV6PLBNezzoXa5+e8TMaxpG2M+IeniENhHQInSJTt0xPr3ZB/4xTxPjDpjDJJk
RFYGA44QpgYKOFZmg4SGVxJ799EO9u0L7ug/JuDODkEM4H22VPxnMtG2vHO61jyp+ege+46SGOGe
PBPtH20/hk8ieUeksqfaZ2pMmc8Eq02zm6AvQEovFdqY6z14QPvEKsyrE5PKFAxEATxYpDbbcsV9
BvVIepddxdywW6dd5CFoy3ExNOrWmbWjOyAiUDQXe37PWBl6B2eDedQprDYfgEBk4YjkIa73bUux
WgkAl+tzGMHzqzJbYY5GdcmM/e+ikeIBBWMIbqCyjywm/FL+MOfKF9l+xWCNhbHdT4E22lX6QZA4
SQa8eiLe8X7rbC4RSRNSY1S8L2jLdpXiSyB6CL4/u7p5z+pJl1QyX97B54EdNjq95B2DZdgbkYlQ
msaMtRqbwh5B2Wc4JCWJOQhxOBmmm1KArIpNSrEL5mlMDuQRyB253xrUC0xrWL/ywEksZI4LbGXW
xaThQZWRqm3UMRusePfnTTCCJC718sDQgSyoP2DgJYHr62X7S8GNiippQFNkGljQ45e7wO9X0vc+
4yWAd0EHvGutu8zHKVAI3mWTuYinlH1Xr94EswJZrfmZcbsHnV7bVZB+bRr09pxoIojA3i4J54uQ
QfUGXbzaWXXdmcQAm5+N8vxuuEqOZon4KdWhfjGPgGPfOOsPXBETk8lsV1clrm+3fAaP+u+IZwQv
udO9x+Klrk0F+SLwhq9F6qYRQqUi9DmRLrN8kLQIJgmZ9IXBjWGXS4028y2zyIuHkPSfH6oq7r2v
hCV3JvYawKqjw8LbOSgE4/rWCZ+5WRio/3qCYYiqHbHysxZQMhxg+U+EKyyUiD+lfqn/ILOCzNXO
yOTWjx5wHHrzRLkOdqKygJrJsE21alXSBcOTZMdC0ukqylT4dPO95QnlgeRSSv/MtGJ4rkyRe8zt
YtK2UBx8HCOFcrysRNyE4IU8jebizRQv7gKsGkkd0sfUnj+IfkY38pWGTD91q2odFo+BKjUvCn43
N11hImQYEBwpYrpOLnFFhB64pmSs1YqI+iTVLAYD5WbypaSvYUl/lkNOvQ4wz7QaAO+eBg/BCX+/
lbuWQZkbo65tw/gCyLPOnAj273KpqbSe4bGhkkd3txPnWi6WLbbBKe7B5iN3D8vkSjFAPjEZt2i6
x6ZCpY+DmooP8JX1xkK7Eee8w3ZPDvtzHJwq420ARWAK1VLl1jonDnAjlGk/WK4IEROlH0kYCB9H
wJCAEXchql4kcguu8tEs54Umkmi7hQxVqGwo1ldRbYltqD82vsDweD6hL6vgToq2fZdGunkfDAoi
xv7wrEe4jTcrplDnv7oSqIcdjmzxZtrC/R0DiQdgrmYh8wK3m/WHk2d+jspPuiqtDg0UO0ZA0UjR
dbMDJZXi8Obtvhumln2KxhVE60YjtoTDLKpQie5MtpA35ZPX5bB1QRkovV8v8dGHk9tA3xLS4kCZ
nDIJDd5C9zbxZ7qaCXJsSjBCc2lFWIEzV1gDXg3NBzV+8we7wn98TIhFDQpAbs3WXw4RqeNVljH6
9IGVF7AIQrWLd4eNC+xi6pvnw9XweKLAfnBZexfu34zOsfWKLAyeKVtETzrO0AWNQCTx2bHTTKRz
Kobjm5ZarqoyhbnC9XMyN4LqOr2B8UNGMMnszNt6jIlYSQtNZW/SI+YasbgKf9maC1eYB7ai9nNT
4YUG6Ha93tAPAm95w2tMJR0P1hy9Vx6xhUQQdWOhmd9WHjEOx0qWKPK5tab3f+/YvSo++toY/+6U
0cwmzIU7m5t2TSUxoEzIDv0be1wfNafF6GhX1j1hvFVeA9PngDHDdLLWPazBgFtDex1hKWQqf7fs
XBGwXFL1MAi1mgsq81TKAV0P5MBY/6hLvgEZ/AVup+mqxOWtDP3KBhQrdqq2bmQJJYfNV6Vw9ANf
hJtl/wDGsbK3XvXoen1tRFGhzWteIotjho+W3VSMJBaoJPF65rMc3+g0N2/l+rJt445C37pzBWBQ
BBHtLUDpMOUnNjPxfc5vQWYhyYk8BPfv9wqS5Pwn72Yn29xlJe2ffOZG7Qi3m1b/pntwjbA7gfi4
Qnm+YZfwJPEjfFkg1eqjIqW8kL5ZrgPklvrJdaILYMOUJZT73RqV+iqd/mZ2mgbSZZGyt5kXu0Li
nCchi69F/i3uTaX5bmk+oaaJBn4pl7myEx6GLnfIoaPLubAbI52kK6zNyI/3/Qaz8O4I0K5Ra0QR
2zC7zLcNW78hdZ62qhOhzYNkzE2kXLCjhH1YzGw2e86Y3tWCPKc2qnimTl+LQvGCvdxyBZ9/lmXY
JU/q6AZvG3TcVQTYPs0E+uiecnVZ+SLd1yd+NW8WYLvI6OTcLKg5YxWC0px2Uq2MNa+doCXVl6N1
1cOeC4p7AFDr2JFmj9SsXhumtuVzKQH149OgwUS5UxpINXUXXjfgwG3ilpoYOES5/IKEszpPHcZA
/9t0Vov9qBoZIOwOi0YtpZjxdTgTpjwFUNHt5Uz6vqEaaGD9UETi/Y+1KBOXG956OBiJ8FPj9VTF
crfpTL7f+aqvUYPiTnOStIyhtWL7WFdf1Sc4bBZy5zWSnKEwe7hbuvtqI4QV7cLH2KqMKsYyB+YA
3C2CMryNTF5ZisgOHqg5rAVWe+aoVjs/hWYzVtiGAj+nNG3IC3aalZ0NQSgmlc5GVSSpKybV6iYm
/D7FSXIlZGIix40kidnAnHkyId+8+iPwkPicgGOYrI3Oiaq91CR/8LYkNRC2cEMlbYmfyFy1OtQk
eVeyL+6nHbF4mrRa1E/IDn2YrAi2jDqSMuIhIwoWNau8pVQGwunXnBwixTRZVTRMfCdJ1qct9GtO
+8xQCwcpE9NW8bKYuDFvRXpSoXcCM8eS7aQzxZtwzNZ9RyB/LXu599Kj18IeqpswmvcpRk2e8E4U
ZBCEEOHFjVX5tjyvAThQqDWFdxXH0ChEcdQ4oIdqExbKX6xhPEkr743oyysgI7j2JSWRkV6hOfry
U3yyirFnwNoQihi+td7zldbr/DjrrnBsWYRiXh9L6l0QCXgnDUfpfZoiFZ2Q+rqGctYkxp7/xTXb
6cf4TPVNqrQdaTLwgn/5Y1N+w9O4XicgWitGB5Cou+tdNkm4RUUw3638vldl5dBU1FumZgwZL+8o
w3WndXdKCIO68izswZFUJX9QcaFkkXBzFzJCOCnXnQAX9QzplUGlCS8mmtdwISaOPxBj/cMsqmHv
V8FZ7QTiSFZlXFJHQdOpafxzWbXur+MY7yrYDfXCoq6+/gNeSOtLzYp32lFUtvlm5I83luJ/ZcIp
0MWeUIaq77RxyKfUNpNn0+HOoOVt5wM1Q/ru6kYHi35lrhYtxZDZhnsWwlQLwWX0jymfyM6B/iOm
q0GEcXiaqnJ4xVtqPAZ219McNU8MnCyy3DOErzibvXffkAXP3YEibDQKdWZzlMUUp3lQidxVk30a
rvYym7hqDSKv9kEV82QhEWFxT07Sbe3TnON2ZyQU1WQ6egs6j8OGWadogA49DvzAZODFjYoLEmWA
mLAJYxG4btgUtNBm2iI7RgCNXZpKyNCvEb55XBFjxMF7MeFIwdmOP3dLHt6WE+XASFFsZYg+brpr
CKcQ5xd3bgEDnME2dBLdt5V7qcSkDpKoRxRF1aqWrFqHu1pSPoIbkWlQuKPSlNrFoHgulEyn0spB
TSRa6UX6KnE1T4Esja4/R/opbEhf1V5efquh3CfFcv0WGgoZqUiyWGE7BuXlSJeEhJwnE2+oeB2S
mUGQIjfbfedU0iKano70HfAbAkv75KAze6bRY77TvFNn3/ZK/iYqZ3R0317bnkHZCwhB3CO2X7uR
ec9AKbUHv/veHsOpqbbDC9UM06ebCL/Z58CvnkKdu2ulTrN2mvpRVQj8OK/OS8s2g7oeCYpexuSQ
do1TIfpkgB+4FaJdnsbbLuwJGGfIlSsxmI8gyga/CEPCHjmUuHCuLLKmJNJQrp0XSPgelPmHW5i0
Md8MnkRsmMJ+nFULAZV6KqZCYz2Tnio/VzgfF5nR3NxYKtndVSyV32HpF0O34/ZP8jlG1T/ZjrBG
Csvi6nDQz39k6iP3cdrKkcFbUlVgL7DaNBgqUNwcwRwCRFrvp7a1+vKty+Tq0KOHyNr3oiVo51ih
HjTdSf1PEZn0AGl0kO3hL0cQglJB0Hl2BW9P85lsc/5RO6a+aPejmd0JFke/S/s9samybfShOCqI
TWxJ3UyU8lrjKX1hTMEq/pYP72YzqeruzQDqDXa6Kr1FH0isIQWD1RHx2p8mbekSjKaW9usfHGyC
yRJ0hGoz60NWia0gAdsJCu/Sy49ITPgWxZvq7dUFEYrLeISJbxDcnG+qQ4a2/Q29spEon5Gg1HBR
twrC3t1+SbF9ARW3c/hz3WVRZ94LkWKTULeeAES6vhZLLKWq5reW0lTgOPjJSCYewc0RMDxFUXDr
8XyLq4mr8EcgKgGT7tEAKX+G7muewTXx+S0Pck1auMHHGJQaZeeeDiYcSjffS+q5WTljXupNDTsS
tplpFpFAXDbZCMMKkMkwW2m0/dZLsNwYd/rUPXfrfQlFDF1uWNCz1UAgsjiKPlb2fdJkyXDQlhlb
771VCBjRI+lwmjKmytsyhMtnUGotZWkDCG6NCJsEnXsrdB/+YNbexEqv/cf6a74Z1nqSHYGky7yi
sg6fwmANuZ5CJPcKj4tnHTdHA3nZsZYwIx13j+Q0/2hJ0yxZmH9fyf9EDt4yzIJyb9QVw2ORntHp
QsGHTY2ED5mM1RefzrDoNVg/c2ql1rv87lgzPrkUL9Q3ySrM79MRK7noCGEVypu8uUxV2aJG+En4
OseSbNweOu9fJEgZ3J6GrMuX49xBTa2jeEzg42MVcgPH4wFVT8IXbeN1jyEoWHZ5vdoB3A+iY3/0
p959b+pt+9dUjNC6GQdyOhqH9WU9nPJ1QObU9QMQwFUbuqm5/qMkpbf1Qw7wS5YPktAhoJuASSGb
ofdZhDW1T79ilReqAu5wwR9HBprJ/G/mxGQpCevNeo4iChcC6L2DFpzAJMAeqUJlXSz9r0aqXhyE
tfy87DUv1K/+OM1bgo7iDVf5GFjfcV37USX/JVnYORtMLGtZdh3vQSFeTaJZ1jyf2gzHCM6BPSDS
q+aqzZfXyJwIb41S8S0BY+kNlsaLWuSmU4mVOnp52OWqPCEp2xCKdPrHV9vA3uWzHMOQ4K2lzasi
e4Ig12zABAF+igU3QLX3anywaAtC8DZEY/tRHSN8diuqLSeV6oar2KjKSiAdGodLWTUcoA984r8d
aa/z6xFAfo/kKKPzlTBSynVhJYm2NUhNP+VwPX9Wh9RG/EHijIyVYMz+crro9/lmrz4A4lGTokdb
EMCd9w8QDFv2hqKlq7puhKWEnvCf+7Jx1fzzpgqCGKCsbCp3/eO0fD4tk8otmWL+WrNuw9ALMV13
qtv4Mk22VstfVmQOspEP1LQlukEM8kcICjWdG1LZpEKRQygnx/M742nbeuhWcV82KQzCEq8O5Raj
yQW62sNJbtap1puYaehFomgULoH3+ifZdIvC52JcVCkThFnYxeOhmChkBzLNmzZ+MYzsCEvoUavP
4w+AGlsd5y4evCR8R9Z3j+DssoYrBc5TRPENJLV9Z9gMQYyoJFhBmuLs/lx155EaG+u6weXdOZ+l
j6dUpgPeqpPElmoNBFQpsjteB/r4/lLyHq1C8iRmky3gNe6+7FtK5AUzbhZTJrUmIcwLEk8452Wu
jHLUpp18SxpbB4ihISgAgWMvZsDNblhnhDxa1/A5/oYnIc52a/c1STH0VQqNGZJ962ybXttpiO32
byOkfpLMpbNhxieN9iv8hlgFqDC3qh7UuAMlD46vO0RqoxUSURo4mMIRPUjXtAmRWi/vkFi2dxk2
DlDtHC49/zXjqoVfHtBh6DAiC+7XZG8SyTEvOgLbuexGqteCTSH3O8oQ3BJPAXfmPI03S4K517Kp
P/QatlIWvi+37idg9pQsHSl7cV89r6FjxiT5j0tfMtdh/laXkzwKKqYkYh3nOIF1Pc9itKeux3Tu
6nZkTnhsKu5NDnVAkfMdDTyl4QhdRZjtRRmVIheDuzsqFlfju+dZ1lb5lPmKVkIFrlT4GuXekxFs
vQNrtWR4mjBs5AM3JLH2XzAHhL02XTsq0U3+ZlKrgH3+Fuc/KxNIxoUKCsRrJZVHI/8RNVN1qO4q
QZjOOotmsZWT/OqUqAvw6XecQtG9jxyqkRrEDjTrKf/SzzLFWP2Y/ZQE29bTFfdLWNy8/cgN9KFH
onIM1Tt8cO0KOK9avXIDt9vmuhJn61uMmkoOikXWcJ2oV5DevdR7Qw6Cy3rAQhwMiQLw9I49avwf
Qu4uRZq6EO8SX+P/6iL3D4HysTRDp8XCQbJNh2IXtDpcPFUsjJnkaEz2TrDYEBHtEwr2/syK/vB+
G/kxYpB6PzRkFcRSOjQ3PImi6fspC16XX759go1wCxu6epknwklanuGg/Hp0HI9C/VlZiyOQmopx
oa5SQnpSx+xhyQ3K9qlgVh777eg4uHL0u8r/sMlxOSounpe7FMWCZZBVQhr9YBJyFRDdkkePNdG3
z64+YN48uZvf3FPtoxfPoZoq6vyGzX+4Uc0cKinKxuCLqOcrU4ksdIUCPabZRhc8GlcI+4/RFzPz
WKMyElU66LfuD+zCXl1AqZLz3Lu0k6CFYXdk5Gh/AbDqaJWKillBvvV9iPTdvDIjRM/tzvQfmmy5
oCjACYyt+GJevCSvZWxK/AOrVsU6bj8kZgbe15eunmSMHcDTuazBHJSBusIc2XE94vZH5w2V+HYM
pYaXubKA+biPcfdJC8XR1wqoO3N/JuHv5injiaV8OVh1R1OHqrHhzWQdy5J8Vk41xL5cAEn4Ag/d
yV/eqCfN6Ns42P+WwCiRRMkyCH91Qi/rDxSX6LJIRYKhC5+ndY9NXlNhMfMgIdLnSFz4cFdpHFgj
LvgIlcgVNQWTFjo6vp5Tf4uDtJSMOrkUyI/+HuUA0pqQzA4jQIIsx95OUzbrrSka2XiYGO9LgYHN
eEGgvQ0NmSu+3pmrXENGq820jgGIVWcqh28ZJKxgfuS/CLJ5oW/NXJfWHBeo8gg9vd2Yh3ZTKmmi
E92VSzVkmh7Uf6smT3Gj2DYvWOITGDvzpvy/L7dfnU5Uc38eMKU1liaX1/0hXivP+qxNdtnm1S+8
fco1SpjB4I17nABzHYF40rwpCUZH1EqT9nBKqyFbzqcnS/Udypst9GYuU/cnB150grvC5gOv1x/Q
O/uY5TbKjKBim1Syke8gYTNNnJSPEctlh3hAeBLV829/kA5kKICeEYNd40ipSNoEsG5/TOiBi3KV
5IB49apH7oDWjnM+IZD/MvUQKWwbQuakVfm7SSlOEwnvmORdArQ/fgH9YPp1rXSn2KcnMUWGBGgs
6BSQhFJeumBkegvz3OoPL4KCUnWdn01kcUn7Xao4LEPzcm9w9om3x/JWJjvngZl/hj0PeIEqcTUa
wL+Qd8XNY+OPC2mokUXgVIcWBZizZzWx9HWlyNVmHeiTGpn4YUD6Z2a9oXKb8OB66IvNLFhwPikT
OM9l3SaFP3RsgiEQwS8ie1n4z89gECLv2TfMdhaqPhPuCYfFpvV8yGBRGHX1weohUOo7bNJUgQtb
efU2Yp8AQYbE+nTiP70N/Oz+ra6xjH7+v5ZK3NGSL2VlEeaZ4A0RCnkXCCJuQQZTJTJjlj718wAT
f+vnvnqGmADq5GZFRaa/HGzaXUbGvCZYCYNr+47LFdUpTjbuJ4+qRmW+R5tCF+3NZyJgwSFQaWyC
A5dZH+XrZIuY/vtEwsyjrWACyoHOp+SNVmZoPHjPGK5u7yM0jKMnPPxMTdzvzeo/5NxUFgkiWQZI
fd3/ADznHynUvqtXZ4dMWIY7tee473FIdn9N2cSx4HlzZKcchJBpYzBUfpOJbYIkpeg3TYkPhlme
oTGFdo8dQ1SCZdzgCfmc55HZXkAsUSt8pTxbCf8MBqqp6jiYUMfi2XMQiO/p/LSDaQJzHPORVo6U
wRkcpNolkMEL2eRpIcRCXkpOM9zlufhPaV3NByaNdLcXUleHTcIrzPeG57JFTgcgOx7zIbSeJjo+
YwGhzyLMURzH5fkcT8OWuDsIQxkcVChrD7oq3ynlWkML9SNxvKn1uH6fvz+PM1WuKALTBlSXBEg9
zfqaK1Ytm8tDgNM1ttV7sVcpWX2lUTCvPMLfbIiX4e9jV2BGjd/tFnE2cPy1H6h4JTius9309GJ7
7WrnYku1nq71PpmQ3dcVzmvzOd/QAa91nuVl95THQOqWiIRqSMwzI5YsIOm13ueZC+8iYHaS7y9w
/T4PrY+lREzd15sM74/1hzyn3L257Eh+UJIdhJilSAyB6w/IKj2Xl8KyNB2NsGoo9sfgX1ril8bI
RJS0G2xw0AxcoIkUqGF7sEom5HwsudG8up4xQGnbQtAQsuJvnkxv/S0j2OapWnJxu6+mzofZNJrd
8qYRnJdumidXSoAAADqR6a2XNhX8thfezyssGfLomJNIVYJY1fFpBFcNnY0CwdMyMv7GKqbgmWhR
mulLgKyrmceF0ylYIU7E/AJTf2E8EueCGaom9mE4sFe860xY5Tabc0TPBxR/pWo3TnfaPBh9iGrg
7X2wKiGjzFKNeThzflEdrnrmslVj4CCGTg/QAZsfTxE6mFmsj8MElhRTcxHBblwHesBSDDi85EFR
fm0Sp19xmlCTA16BkoGUrUOlE8Pebdv1cYJH90copL4+K2Vz7l+utRZuzyPAMl/Mi+/mGU3kuyWv
UZN+wrskQEJNV/jLDdQZ9RbXkQ1Vxa/44sGBJjLh71k64rnI+xURTCfm46z08OEsWbjfGE+ZnfYf
LJ5BW1QYaqP5lqwtA96oz0KwSRsc2GUmPYcg+NYboeSJc3Y3Jpaw4DTY6L2D8n2rAbMPbAziwWYm
1wCeBICoxuNu3M1Cgikh0vZigolBsSwfwM2RqHLEkVIDvi7NJZOtjB5jVmYsuXc7WiDQn8mieP/o
NAhBa3kJgfG1JSlNfsyFC/2zXk89BbsL3rHaEbLNJ5dppQtGHlw0GV32aE7ETLi2fdekRwO/jukL
v5kbVUlRYXRLf/3GvaEHZbDRz06kJLe6YrL1cmsn4qKTQ7jwMO90wmBtuC1hyek2MFlfQsTOsxr8
nYIrlJ3nN39nqyv83qylSPNMn+R6/Mx/xBgt4nNgSnfUdHeLzr/zhe11moJ1280g/u1Z+0l0p8/B
EevaJROjj3zmYefC+/D/qV/As+EnE18xTcRO+W9WCCy0iUKRRL1dNzJroEjkTcSVDW2/htFYHCJC
EEkLfBm6yPy7GmscGPqQ4+1/7sN1vyahLdy89mnRq75gepIiUl7fVxNpM9RgXoWg4B35fmGEpFiZ
TaYkKdyoIlxCMvlsp0GzslA6FzxcCJS1EV/wwBDpDrRbTiyB1R9Kh0WYb5VLvRazjdG30IHl4jvw
mGGJSu6g0u5UEBFUg2Tw271OYjkCAOIl7OuayYdZybwvVdkqCT5DLmOGu6AQ3nKI5KTzvl3aSCPe
dsNLfQhEUnF8bVAJ8ws+Kx7Oaj2REPDH+8DZ2wKZ4kYEIDH088Utp/ATNQa8u9kGrhqJkZBDjXu5
pMJg2R3hjvun/BQ7ymmfL6cvMYM+T5K8yJemJbFrsamjgKRwrB87LefagXAkZaBICHMHmQxemGHu
SscxuebweBC9vYi2sjGJkjpYQbSnyG2SHbst6ZtLuLmc1OJecTsSpEBap42b1QkRWuxgiNFN5ieI
K+B6bDisMxbDw6pbgN4fsb8cqIM+y0wifgO4aDxjgUUXZ6EnplNkQZo4ApCRYojlbVHm3mc544zi
4I49Myynk1cVp29td37hFQjlfCkor9DYTp/PtadL4cfgqzVWPANfqJ353h7H+1LNFrpL8DDOa95y
3L7vYuFtok1qywua8BG/HV0307WEu0w8czg5EVlGZFMaO0BTHXrPTJS27C9bQyYixbPjp51w0Zv0
g/RyYtg+FX4zqjltY/MnP/N17EYiOVFGZeFk2v/XZyCC0Xbu1yZgFSY1rTRftLunHzAHmAkaNbhR
l8yNkz/e2SE2r4aX53/aERA1cY7fbgIZkS7pLcn5LCAwejIEgE4gzVOtMaELtbLZnlnpdJEt5gfi
83u2CLGBbdKrKwp5UU5kV9LGauLx+kbYjEE/rJXLl9sheEyxjsnJ3u+uLkXjjbdKmlwbBrCHdO4R
qqz6Q32QdYvXnpXuvfQBchiYNFOY7BuuJhKIURjsxVQQkjH0mMby3d4l49wcMb7qQLkrrPVir9mG
+M5mN5V7l1HTi/8KzkuQZIrx29+jHfk2lonTN8/pdRHWxg/Z8tXaUFk8MpIjZoRG+cwUzoXMlymJ
bJJDaVa5yrCg4n0HaWaSUeE6Rh6JQb/ObOcWkq4UjPtap5bhpZuzVVJt7oeDDG5ZuFVungAsHCcQ
v80KIJJtBmVbhzEeA9ylUk45iXPBjk5acd373fVQXfhY5vbhTmTlq3GDUOwJxnGHMunPVP1Pkcrj
TBLUU4Uxmwlm16QW+Q4Pn0VA+dgrvSvJjakobvAiT7zBnTYJ6odNk3eEi2i6X792rU1w7iRZ93TW
ct5s7+gknMWFC0YFSdjt1IWOkgSBe5hnj2DlDnG88hgJ8ngpH0WOPiJeAORRlIr6LPLpNQoRnrlU
apvObb6nnu2mcy2P4wzFohBVVuBq9OwLlbMsYIixab4GAAMfR/5SxaKcD8uPQCmB4wTOrO3OIu1F
zl7+1yWkxYKs2aBrLdJafh8aAQbUlh0nse9xjhD2w8jgtXZsHAHDUbX9HhEyO3ilSskytbTYcBkG
182rqv0yW8/QvpC29ozl2NVQ7f/F6dW0D0zQZuIu1KKv42AA30UiLCYeoTQgGPY1S0LKYAoJRyuB
czZbJhBKkAwBVjMGIzIYSKoMuUJe1d20jJEWYBfgHJpVGb0KZ1YQxXetbZhp4s5rBtdenA1zMZUo
wcm4MF3u4C7f23fZBjqoqlh0TQIIb08RLIAq5rHFI5h1dhX4lNYGADlRIC4SzImGyU3s/CIuPuq0
1ofBx92YshZoDRwaze3iluGvdI5lHSq1iKJIJeOHCdmdsJAxnt6uubdqD53+aOR0IBnYssltDHoe
0xmnRfW5m3Mk7AzTWpF5BxCOdd/dn+ytCMuUfYzJJ1pfRUYh/F6ydHorX0h6zGJkf+8yomv4G0NX
fMmRkbB2NbXbV5e2+tjyrh/ImGp1MAkLRJUQbfWfswe2PsCDTxF5zGUVqdd1OsOHSFjWGryNnLjL
3HiY658PDRTIT0vUg1I+iradSoGUguVJUn80/A9vKn7Mcuk1tDjPkXRo1i0LgV8pkkB9MQWuxgcW
JTR9Sht0Ta79NGPc7iPUHRr95zISsOwDIWwvHHZyp9ab70ohMbaBP8n+EohE6FaBHtv5/Ut/x9D1
+4wFyPKQ542RIgXzKzfgRW33auwtD3pizSfpkhFgLHGIGUskr3wbQaqEJxHKWqHWZJRlu+cKKaoP
Ozmwe9fQxR0dSDmU+hOe8z7NaAKy2mnj8Nbcysme1iTQ7dFZ9GMdjqs2+y7dc+fwo5ubT/1H7ahW
B1+Em5SV5oAyPMT7TFhsufcTLKj3cwYJ02bAEYs4t6RuW49fiwHTLvwBm3OSo0ZV+3+TFvOSPRrT
ZwxJHd1FD2r993voBZzH4V/BTWhRsLWIBKLu8RzAZ4XOGiq0CMHkMeMh5TVzM8FuaA15Leykvl6w
/dpg+wRjFII1plaJq7kVN9flCeYzUFyMpG/8Jigp+QUVJdIYrG76fHKaUqymyvs/e44Yxnoml7No
chytnm60D5iE5E6uxaVyrF+DpZRlX6Nc7lAOldv/U6zXeKv/ug+9FVP/I+SVYYD3z2ATYsT/Xqjn
94Sc8MA6M94ligpVkmCecEr5+o+2s8iRUwA0WFyz12eVqRIWXvmDtwRIn1V8wXVE1agOEEJpvo/P
DJqoUuRisSiwyIqbrw0iMl3fgxPyUwD9mQSgoYwKiW2HMY4QJHvd+OjCxY9KXAx8eU8A19q7uZVK
8sJDpvyiObjayh4Wc/Pni7kQyFdZLvBorgTz+kvY78KJkFvAu89qefI/aDlp043i0LvTo7fNZGl8
MrV6K97wbnkUyGVqg+GhyqdQAT5E/jCJjKq6wDVH/8WE1c83xJvgSbur/d4HLc9IpfM2wmdY+iVf
8fV5JgvVxHsJ48rW6YM3hzR6TGc43j1yzNw0aMwh7Vh9JSEFArPMEbDZYCFFkZ5AtHCxMwwxaZqV
iEXed930CtuCoam63Lv18Xudq+7ZV5ArezHynqKRDRhRx8Que2+gQXliFNmcGDDqos/ST2IL141U
Y61MNUbQweBDfPH5XuiZXWJ2607vJ36mh4ZOuYnj4juSZtJ4IUJXW6nFqS5Rs/cM0KcouxijDwx/
WdyGuHTKnC6QqRpV/laynmjBhl67fq5NBKbtxIEt1hX1Nx/dLREeCYaf+uNG2ef/6RIuRAsuo+6t
WZzPFREvoBzM2NPIC2Sev9o+jrt+/ETcPwxHAP5u75nHky1Gcj3Rxb1jZZr7hSOBl8ExU9OWwMXm
ygGyrOhjvi7H1Horv4fD0Th2XIES68i/f2gZpfMV9LbxiYsC7d0BCKbSzIr5gifoABA8pTlRDtac
GmEwpfxyISomyo72aTN/jBdrX+VfywwckxDJ/kEvn9B7syFN7C4sTlH9pGsl3Rqvcmsrwrld+Osy
iAk80NdK4kOkIr8/NpUzBuqj6FL7C7k+c9Kx5qGFC6h4Hl0ZrKCfzOIdR+QER+6tGE+AMF2c7yxB
lFaAJRdROWIvv0uToelCM39PVH/RzOEpB3PwD6+OXfwYSOl9jjNNScMrmx2UNpiQIvM3OfBGLs9V
vj0+pv+V7QJC4gl3tH2SKuysnF7oDNpC/IXR+C8AhCmksujh17gZp/VlfTxQbRVXe1PPM1gaaEva
cnnS26xnTKv/zgJ3UsUFPpUq6xhWV2JAUg049BVLK1H/pwQqe4RxDHdvGatp5KlL/8/V5cwsvsis
i6vJTBl0C0wtFL6bvwNtXFEdoTHWyNKduLr4qtO1Z8+78mNzFhWrqin/RsiWoQ7JQxBcflLwr7kK
Whie1Mk5pmZv+gL0Dua9LS/8nxCz/7kvKxblGlElK8+4aSOd9+g71zONYQCVIYdwK2AdWcTK3X4L
AlQFyNsstZNSo4pNCKszYpET3R0td1/6p9Hu9PhyroBLpb72tRjVcewIxNC1O3ieTkcfPqjwxs5S
VQPekWA59sx7AwfWr2g9VV0QFRkNcRf17k81Q9/QxmmfwXapNtFIA11Les6TG11fRLpRjfdaTtTZ
IPIbc6eWBRthNVl7Xye+xuBarWXoz0Yq7mEoOCaaJUcxvhZXvAn+O1OjFBNuVQ4+usgSnjsnVyfX
Vk4SN6Cw62CGxWpJLPj26h5yP1uRedLWL5Adv6n1CVNYufFc+SqsKQyuQA75BGRUDE6HURbAVhp9
Xk43Wtl7Ej6Um0H3o1VEoXxD3IRU8zSUMsm7+0UdtKkJQMxDMKLk4l/JBJW7eNGIn9Pkarc6zuJ8
IGIj8o1+EsYitPB+LE2QUmxYJOq9XRncw32rMTFtYaMFGkPf19ZTlhDF2Higkl+jLZkcxAdAaEte
LLQsAQvP+DK9JFcn56mtOipjGs1mzr0ZH2N1ndiMvsbXDhJMghVugDVgRMi7pAui8FpBZ2ZzREd6
CNXusZuZtHsakaYgxgGa/KOPGntSNTwdg0yiM+Qo8GuCnVfBCohGEhWlZSbayFNAbH8dUGRgWiak
jJfaL0kE52YmU/+BmUjmYqzLVmwBgJJk5iRjRjZxldVhl0WbY9QZEauPgpFhyHAQQZWHF/2/AVpu
TZnLO8/zm+UAgzTevedIahNEZoDltD+OcB9VxtpehQEQmofyf9LryGhpQL3laZGYNEQ4uf5mAZ62
m4BzgKnqgBAvNJN4ctvKOSpc4U9hQbTrSLDL5PGjkSPdrCTa5RlGm0uMMkGa3QXWsLSrigENe5rS
VroavuNkPsWy+aJkf+muN1rKSfhCiEF9DAuSc7XgCb8wyUBQiXv+iPH0yDhCg6hU+Muyniheab7j
v+//qfC0wE8+wFD0dZZ/c37/3PSyAyDpniWPzTtKY8lFOow+GlPaQ03GwE310pEm1JHlg3Ahahds
4+p1rHxKTEBmFJSv+OMW9TFJYaxIio287MAXZxYq6dJ5vXgzPfzIs3c0RiGcTDlo9uaeln0vLtFl
QPhH611wPnz3mirkW3miFz1p6ALRNYMZsfv6wfN0kBSxRtKMT31UG9TCw3Eh87Fj2yITcLjShnpB
1umDTcrpXvDgFA1UAKAjqYML4XMN47ucBM6ujSXVZ85ZOp/0RuRWDAFT+LfubbfG6MuHPjI5cVbe
MK/YHFWBkXC3DSQGwbaSQjQHz+SrMNYnkNZrnyi00ekbp82QbYkRhAWcxPFeazabHGnBmvdRPG0T
hcgJYSbhZ5/yMu2K1Mvh7VdBCI/G1i2U7+Zlu6gdGffPzhQkLe5SK6wWJFqRkpmm99ApaplU95iS
J22DNUq3EXzJytpcFZJbqwQtKHyT4E5t5N5S8FtqBHXsFlgzwyTUQJI49PC2gmANGbrS90z71pTx
Lm3KJTIZrarGM7H561qoINHsHa5OcUi8gO0RFj/Bj8Z7bKk4u3l7ThAjWOFxhNLOR4tYsnQs0Vr5
XsmWTKZL3MYnVmYj2L9N5h7p+3zPbGm+aJYkDy5mkzlIY2zuMjY61+zJYXD31+fL2opNNnSBsQFV
4+P8YZks12QxVqW3Wgwz2uz2w5NzY1RK3lUIUZt3ar/MMfY8WYKs/HrFCpYx9azIHSosF9Tv7zHS
Vyo9QqK9qd1EF0VHIiBXYv4bPoJ+6aYhDqFxmNk9IAbYwLEk74+GYpOKKqdbqjidyDlejL+FCm0e
NhgEQdDEgqVJodSnx1T+R9kZu7+D/V7yzFqhJm8iMvqi3Re1LsVWsiZBQz+cMYw13AIKCRv0TUu2
PA5PZxuSmIxYEZQjX57SJwVN/bMP0K894QWpVgFGyZjt2aMjBXCsuEDRZQMPcfYrKLMno3zAPdON
FXZK6JKsbAZiie0OtP8Jxt/wFU0J+SjiZrEAb89PTD8aHlyiUqvgxbiSsotG2WZqBJqeoxg34QxU
w7I4lqoDI7egwiTaVMKF50V0yXBUAspQzCFF6paFS1oQbzisOzB+B2WIUAVuODEu9z6YJ1BqGk2e
UTeHXY7XGM6l6Ndc4eKsyJjeTiXUtGourDMwiIJEMjUudJPr1B5Ze56NDMLVwFwhU0RcJA06r0oz
Ts+44o9DDlRkJCuj5ZGZeZbucPZqgNLFLzjJ/92OtVt7GOnzp7eT1G4jNWdmZJ4CGbiggyRNhFgl
BJYtXoMLB0P9IPc/64XbhZPmE88nfik+gCfttPY+3PZAtcX4AnNjHR+xPbtWTeIw5Nc5FGYqIXPn
GUKJVRN6ZaGyk4v1mlVnYEJRI08Vy4+g89WothsR/fuhqUQsVIhj7p08lkJgRVyn1v9RAsddptd9
ptpliwTiPYDg6KGV7dtUv7OhLDN5iqQ35KIQe9xp3dLEfn6jU1VwA3Qj8BmKQ7BQAO60MhV6jymM
zaozN4Po5jlRnzey5f247zj2Apo3pa3jNkG2PxZ9Hl8iSejm9DKabaOaOcVo0hREIGr2sHDTVVXD
gCE0SGVM6gLiiIFUeDt94erLHxiAC+fE4lH2cXN3SkOyYhJ0mVODTT4LIGWO97t9QWXUKcyYYCRI
q414XCDRoDf1Na3WkLkTWelJ2RW6BvSO0PkHEXKOlMLiQMObtHuhaLLljiANg4eCzCzYVzkrDCE9
cewlgJ3qEqMqaEiqLuGdhejZXqXmFwWBaYy+21XFHpDqIfZLIKofm6wc6v67dtRrNybJZ8gZ2GhH
IOwbOcYEnyKQs4mhog8bZlmP04Ww7kj5gkabE0wtKsdNQ4oH9wDFtKv53ZdlxFBJgxywE9NNla2E
Hiu2VvIShX47y/AsWQRIT+/N5QDZOGsTV3M19qwB6+KJgVuTn7ycnBXAg4Duu0Ufw8TNZLuuDBgI
ZcqOJk37URCBz6PijFnhX6qSn1cWCdlDNwzmTvqmC1W/OfDUraah9hJMWQr8CA9KpWsLrDICTFQM
oRpeymF59CX02SKiW6NetcJVIxFrlNmEbVoj0LApYwvF11c/PI1n7iOsDArAuIkYQFkpPRaEAoNj
PF1zXYKDCQldniXwzcR0NQyXnjMemgN2MdFU3FjSIUKhI6uzrz77ceTGj9NG/I0cMyQg20BWI5Iv
6LjJA0PPa6TUJlawS1M9tCgnpUZUD4EmD++6MR3bXXm15BsFYKoHEf0sGIXORhJzo0k0aj55Gzjt
ru0q4SsZu35ByG+TzCYkxbkZfp6nfzn2PF/BvTKywRxf56bp0tOOVOVqyPwph0RWjz6cy1h4CSfL
KAN0PlskS9hWRXfKgWAsdFPikLVC5Xo5DFORgo5Il14wkanV1ZFeA5zvWeihT1CwVLDdlVuckBTN
bG9S1sW4fMCBzFt8/FLHOdsACeZV/70tOo3Ddsyx7/AUy5bYkpdLAjX+FJrH5W6ev8mctoPR8p8/
/ffnMdyeOFJzAUj9ixYf76YdS3OTMSNL6VQJrw2QwBUMxKHPE/J1GE1KzkcgEj1uzTQr36BRDeiv
yDqxtyJvaVKFRNoW1BfX44bltGWh9K8+BVh03c2PiOsT4G5diab1mkrHXBiBya3SAJgFhrAEexQ2
2kcVDA1YHKbkHgRQoq4pvEhnHq/XGcyuFpB7fUFEmYAIuK7tZkNjrEjXSHaBSwRYAQotstLzId84
nO2SPrs113x/2Egs8ceIPkmLcDeokufTDnw26BifFTzsky4USxPzZuwD74DOvG44fTbV2wxHSpig
1Payo8aYkPDqyUW7SxZrPY9LuOHvxbT5G0EA1ZaGJOZj8pICar+5KqeUu1oKi4BbWR9X2aEfaEy2
0IOs6x/+PvF7OBghqelZWn+KTUUMowFKZIRWB+tmUOnDWW46ul9OwpoxZumP2ngeBYQWcoOeCLuf
Q1eAM6vAjSaKPZ2IX3bk4/ISRjI7lWOxCqDSwODi5e6HnrnipbN8bckpuknsCUA0y9BBSFn2BMHs
/jJrtrsQAJ6KDosptbE/jibKivUmgQiSkGDZOmx/yK2iEXfy+XO74IOj+gASDqMmJBW+aguKEC4F
WC2JdLcEhTY+8rVnDb4gMDlzy24wexiYBiaD+PqXDPOUW84rbk0Yn5ygdqMIUoq4vf7JumjKroYd
9CDoFGj/rpvnYdcOSOxWcsJz8uKj2YoTKYzQ/R1Nw9bInpBhLJKQhXkfUx0YrmUmlx+aSvpMNoPZ
B8bXveSNeRLX+/NbaXD0V5fotJc84I/G/wdrti3vwoHWi7JqBjsQViIQ/x5ZRH3+6237VJ0ZrxNe
0FfhQs1j5SqU1dM28AaHZk2ZDh+LV43DuTFgHFKVLIcaWMCBIYuTxzHZ2fhGATp4pFsO82dVZjCd
P9MKkUjhF+FtbawybUXWLYDIcfjR7X4OAhx6L+Jt44fUia/UxDtjBuE7zD9fguDJgrukOE4sBgkh
4tscZ2YNsTtHW9I94VX/YnotWKL/M6I2So5hB1WOwdtyCmviHYb3xkR+gBzUkVKLdEIvMK9Y4DCC
LdvMBSYOQe8QoCXUl6oqfpx81JXOaNMVk0qFrOgmeCivyxxFHCK1GEh8UwkTzpkEm6xWYwEve5kz
k1eZo4sYpumbLcpg4iZFkLXraev3DjdnVt/oCYOAuzGMrnm8gMsxs3PkeO9AoAiutH3cIW3QjVI8
UjJrCN3R7d0mvkV/xgIx4P9/cYUPVDEKTGHq3kZsFpgf8g3Z/7EmWPpU0k7R/keaAsNJeBx990GC
jr/BVYAKZw0wX122s+8W+OR9thWrFRcVgpZdHhSJ/hWEsPWpwJM4wHzVuQLDcxmnxXJpchG++JJn
CfC6+DJLgLkPHqKvSxmorMRjuqHWRTQvebnJtdoKgy/wLdc4UoW3g80lcLE+zxUPupydW3hZEwaR
KoMpzUeAYoB9iDUNRDbtFEl+kQMgqGDfhh64Sla9/IlS0lB3Si7fsQBVoJ3T83wkHg/nJFVy2I+k
jrXQ9UsiEAzy1N/8ltSy6l9tmDUGxoFH0HtxZOYOO1Hze2+KwwuYuX9f++AtepTEIwFDgUypZ5zd
KydBKEBwumvbdEah+wP4bmM+X6CpuEKY9skhx1LI0PRNrFzsYWpKYbVWgIrrrgOak23pkGr+i1zg
kQh30EWapQzAmyRzW458ZeHdb9YIm/sHVx+5Ep7W7vLiADS90kFXhsqW13dppznvY+SWfZ+DgCbO
Ir9oSgjTuz7BdSFuRWlPoIK7ylYL4wTYFeU2xYUVvLlWrK5fGkmGRzBsY9TIxpAv/0KUardHXaJm
/up5zurTtw2e2kQl65L8BwIvwPFpg9jxzp88kbtcvEXgspLraZzpIRIyCpCeof+p9g3/lIYMvSPg
NRG2oCL+t4Xu9TpDdxkRuOeP8x/JS7W0LmFWT+Q/fX+p8YtX89SyGrEGNCmAOO3MkRvhUd8hyuMg
euS71jZ02jH49Nc0LwWz3+wqubylBxI4zdiMSTtlU2uoxhshBofUCdLVSmgFlgKwXUqiKlLLU+gy
drvAOWDPK/MQM+hAWAm04ShbVpO9Q0kv8sHtI/DOUHZJcGE38wzoNAqeM14vWtDkOYXcEZR420M7
LFsAlpYwdQFVMKgSg3bqFGqnd6axQ23oBjMSw6jrB3B8teR6ICyokII5yBlubRQf8+/hbMQq1AxB
Nk7Z4SCyHTVOnwR7mHyfnLPjFZRQtB7RqPkj2KVFm0QT6MSD29lb/pt5amg9IgJqmpL2qFfb7bjk
A8QQCJIXaRuyArPkhnb/qOFS1fUWNE2SOAGDVf7qLfjDWBy5VIUlZ3xmTDOlgdRwhlOHzp5lP92v
0s7YqoARk+menEelReu+2nAMSjToPADcY9SNEJsmUQwh5dHVv3T5mvzE/CguBtZ5kvDGAR1fyUOn
FWYslKOluTLJoGi4MYjXRImAOhhiZnVxUUznbgdwwUOORsO8QndFProntr0cnYW0PYasryXCYFFL
AqYi8P0sR+aY5L+qiXprV/215XhM/BE+3uFltgSSE/nkt3Fr9f/5Qas8CkchgoykhC+dZHVTuV0r
V01g+YUgoe01T9IClLhzKlafClnqMzuQ756xcrnKixV3YQyMGq4FskX63NQiSvhydqk+mn7oXaOj
XzOfCdDRY1cYe/3IQ2QRRww6Tj8rRDcM1IfglBPh26YFYrj/JVj6854DVhVYb0pLQzZb8gwdrAss
Coq43ewWq6LF4kvrMmtPIqyuFlseqEEbpmtzg1pEzVA9t2uUt/szQOfeTGDKDoGKBuGUsf+Lv+Np
s4B/t/v/+KqxfQDxn7Gz6OBx1HrIlHk5LVS/R8l5Sn9EGYfL+cJHIrbs47mxnwBn732FyFv89V9G
5jlBOiFBH87MBys0iGbgO/Oe7eIVyhgtkmzaMyoKhH4XfryczgsHnZFOdmpuFeXIwIZf1BsGFoe/
NLDJRxO+p4fS9DRKHVcNZN4NF5HIANiWPUTSUN+618ErM+RFPAeic7T88jA9EDhf6ZnXRCj1qHjT
RkYLY1jV8clxSunEXk44r8JnUHsOKxeq9XV6zWMyrOGOUfU97k6NzL4MJbcAq/9spkv3XzgeQS98
7Y8o8xlUMFzfd+SFWMNOagGr8e41qPHGsu226sCiCTRFxAdDgr8vxtbOxHeD066r1/iwHn6VCB/4
1Ajr5vYaB+j4GGp5DAc3PfpMfws8hthbT4xk5T1tv5cNysnCWiD/pWMtScbBGKkPPkHUd2d84LF5
WrEm9tRaKrIUoUbQJ1ctZ0wuUn40VKiMsjZks/dyN2F5uuK4e/zsmca3JIn3oZbrfaJZkmNR8CYd
HNOmCKvZiGm9DebQmRMABA8jsczQn7ChmiG6P3Pmln2vXuwipAOimUTvAlsYYTjCbreg/AQ/yUH7
xAM95fFjfxJ4lRsrdYQFNhLGDL4wxhkPGWboBFiMobDlVPJWISxVGHvEMTrn0x9LdAlZbWTOXHHW
kLyOu9lh2wpcZdyHOYWxcMDBMZle4/HA98ul2NoyO0lGYSFfEsA12DXfFVIcjK42JQiHMXsulUVb
RiVQmhT0bL16Emm9d5H2yNm7rlEUXY3LUdMcEyYZtxLmCTyY+1tDKQrzHOmb2SHNyCqRWNLnxxJE
vmwf0cqEldw+1Y3bdIU90YSLnV0KgDHSaw0p7/X4Et2VjjbzGHdRwX5YRi57oo1m0cNRsd2AKWe2
3JwCyPglUIYvA7pPGP1XQDfL+uQTT2lUUeRZGg+Ph3Xf91gFHfkv2SD710v5daDxj2I6dXLyMiVJ
A/vWGLlyqSofuR4Qxxm23hgFCyKHkG6E6R3Zjg5PbNuMpUA4Pqt1QtBaWqT6Ss4xvyDtPPbqeKpM
yQ+Jvbhn2nELDxxm4AiZaqI6wWhweYU/42x8jXniEIxtEBiRK3z4Yf6lfnARcMHfrHw9RMHCZWJH
4lz6ha+PYAxHkfiyStvsQVZ86fdmN03n6By2Qegm1tAa02wzm9m9V89FZeOXQNHO6wzrfUjtaelB
PoHQXDkSofTI0MQn4FO4g5afXWxobyOc69pgqI/SbMjk33sKH/bJlnFfhN3d7nLUi4agnU/DGD9y
Z5MEVaLcmHDNnhf+UshiCYZY8Iprj7W6yrTPipxsgs1O4Ss/Wjf6GZtmqDM7diQS2IzuJAHwmKzy
8mKYuLq+UtA9jpQKDfVRv+MyGhEbOqZ82h5qiujhVEC6P6GY8yRz55siDCygBGgMIYq9hRUHkCa+
kLbVprDpen/NDmGxjROun6x/j/vNmCWNMrHRQYUt7lHwubmiHQoB2LGuHq6WVcl8d51f8BULIb+n
QLTO4chpGei7902lXpVkWX+YnDYWwskM5nCMZS/79AM97xVydU7/GqWUsMBQIEvS1ozHcXdPwk0W
FAXruL6aMBu3R3TCXw+fE7o1A3SnU1wJUyRPlm0lkwX0V1y3Te27TDy4rb5QPAIjGhOer7Y6A10F
wmqAuIFTGd6EQdQHLgVjSqaYephWczLjurQudcxPPpnNj+Q4fuqeu5FC5ER0nnursjSb6HkoUXL0
E9I8pdR37Zy5TuHY+tprjBtmjc290+SbRBbT22rS6y1gbGWkrhfhkD+DDDEAmjhiY/dTOu+0fwW4
alElhC9nmE78+QArcYVbt21j1RcwAj40gKFFicdztj0tPdRUImJ1iup3X2vCgcO8WMEW3KngBmjM
UrBS2uAzZUFR+p5U66W4ZxNfC/7k8oAzmjzLfpLw+S9gv/CBxvZMNu1z3zcIY9rcUD2OtxvAzWyK
+LvGrRjEidqfmVomgi6e4MsztFu8vQePqbMfKksj3W7HZETXay/rDW8jSswUK1Wleasum7pnTmg0
Ky8YzZ5UPJJ3d7bXq1VAP3gtZHctoo/ymYiLA3uTZZwUIjM5+ijkDZk+xhUZX0hjnaArB4EGZP/v
/ytEj7kxgip/5xH/O1LyQuGorpdTnyGiMDEzOyq5fmyvB9BAXEASGOOB2VqD442SHa3ItP56wMVH
r+k+/rTQQXhvvckHT/HcgBob1ruC8PnUJtnE44LvLiLJvfdiWMlJr7Q/Ga1YhscfXSE0XWD7BAFZ
LUETy+p7z1twuDA+/bEBNHhJo1fxmmpEvKv8IopEkayD4kdOHq0gsDwiG+EEqM4uoXvRNO2Aap+X
cTnWBtxjdAgld/WNrtc/86YfZiyNBGwcHvQ56TQDdIGTdV0mB3nH3nuYCFgEVaMTJYfUDiYvUmLO
aCNWx4YmnReO4XkYE3tCkRV4VQ4Gn9J3oipExOpknrMR+tgB1ZxrcbNfX6VxERk+FsVPR7V0QiuC
+J5WEf8UPOymadILMFvp0sIZXZs4YvDmvZLVsLVoSQY8xVW8FR+yJg+J8/KyyA62i7UmRz416OgU
m9OLPSCmvfI393aE0k2qAt/Xk4h0SAYbwOZG6gBaOVvITJ4J6gSIezVxw903strh/LYtgommb7OY
EoLGk6JbeizlaeDWkjjUZRysOst8UXeKczit/sDIW+Y3O0yU9umdgeJHJQaRrADmmbZ3XlDZAgOt
2bOFs2eqZmJo2TwQlaYTYhkK7XxIoTPTmR0dwmIkY40YVdEesULaQttyjSJamyTcrz+87WmKVlU6
n3Hv13KCxwjQwvf0H8F2VBuQ9+PMNwdJ7OL4ed1ucgC6t2KyIuUHW43G+mOM8XLv73uuvyynkAHF
IMtlNQnHYP72da7GOWGuJNoneiUseI1KJxC0y7ItsKhPoZ1bKgqdtcPgYuEli2D4wrTBQwBj/F4A
fVFQnDif7Yljcc5zqTyW+QnDWK+OljQw+tEwznSiqx05VscQgHK0eJ5utQWFyQgY+QbnCax7pv1D
NAI7hjfgHwDr5AJKH88Agyj9zkf8w/NOUny4tuUN/BBK3EdHdxAdVTfxN7/NBxSL+gn0FBaeKQme
56TsLHnciA/SUkMv7A9FKZC8tzKYS29MCmQzNdBhj6TM3F4uHJmoLaMgAsdzjGaTSBSJNXE4davZ
VKHbOQzOvzxo0DQYZ5Mk3sHAXSDWUYiGy7EH/0CsOYNbGpZQPxTqSuanDIa56GjuBvkBjNuNVA6S
/b/GGWLPVz69oHVClNTHKxIDplXisKn5ngk3LK1k+IJghi4DyE8tzC7ab4onOgdzfdKI2azlPBfI
DlhBNff9eEqeKdPIR7EEwuxw2EfKFCA9Ddv27WLwUVowBr+BbmqgjtFjOBi42ay6sVgo9qNbRMu5
VQzCjpyunaEMBkO96ikns17xzmmjWHhyO1PWM95h/ChYW78vO9vcXPdzxPQNuw2FJem3jE5/kXGe
ioBxrOlMiKkNMHGEQ8MmRh242aGbQ1VJZrM7xLt5lhV1qT6qR1a1EdHdystodut+gfX8gPKh4SsI
R6caZ0TFa8hi0BtKeDyyvohDB9QSEQ/rWt4hitwiGFK9nWVXRl+ooAEjFfpmKiXP+aUQvu9wuVnH
BzHG+1IDuk0dCXLikCYmbhokCNJf9NEYg1WeiiuVCcF6VNSZeD7RiGwMxSscLtyVNwjB0SFiEKhs
ZtMYML/EVg+QlPQHBDeRhDCNks0bxkoIpc5wFqKNjDjoBHvRksyJjl9V/DLZ+1TEEZ56/3TSHPzD
xSA9wIVv5+ixt6FxvCBtUOPLDR5QgTqhMPBqLAh81LZk8tKJbUpDAWdlkmffUBbj9Nfik/9tLWzJ
fcFSqru+BHgvzVagnqygleGw6NPt7cMFqrratiAACC7x2yxlMaZTlrfq0+0ifT/Epjb/LJQWU1fQ
05RbZ7i2AjYjRkq4TxQTuPMpbQoVz2FKIWYzqhK+uS0YD2T6a+ctZkLnWdjXvvNGIGabAH6jLYR1
1X3K8RbvJDgDMAiYvz0DJRxM81YvmeiD9ukybC/2+n42Q1LexRXW4Pja19jRAbonntX4CWy9Zyzz
URtHWxIwYRnBqi2A1v9D3ikUk3/uEUps9jfb/W5azmvFELezfBeA5dE3bptBFyD8b2P1vw1gnGBB
Aoh/yRl9ZPvJpW+lEHanNp5zRLNIfEyPHjwj7r5c3EfvIXYmGkgp6ZFGEOOwdtDhU00cfgXiuVZ7
eXv+dTmr2QmzAawbrbibadqBST+ePDmqwB6y8Qs3AhtdUB1wmdRkGW3yAL0UOMfyfg3C0XSBlqSO
UZI2gaJmx4G4BmWv1Dd9vJoDOtCOt9qRfMRZdNz4Jh+j3UpSPe9ba7sTfXnIW8DxmUQ7DxtkeNdL
+6HapmwyfyAUh8g71YgzPpK1gWLWHzEGYZxYAHKDD4VDwGmYg7hlfVQ/ZAnRwqh1R08RtGFILwJI
zT//puof/uy5J89qZ/WMip6ti23yq//VBERebpnnRA3Ir+RSc6lQ2zbtiFjCl9ikvWthFe42swmC
yC0FmemuAWbTqc93QXQvN0/8XxJAC+IJAmGe5onb4P2bdG2WG925oVW2eyACY8cnBOtRii3CKKVZ
6PrUEmA33SZquJq6yI7fFJzLbh/BG189DRtCbwUtcp/LoWFXm1IDPmh55nxs960VlD8AoX9KyOj2
1o5gxpXNbGMW1Z/R6qQUQ/gsvREnRYF+GU1rNIl20+AKIUplT+iCpjtYYIVUCk5NXAcWl847MFTi
hd3NyzhqE2rfiKSl+fbAFSmWrLLTWEGpvG16ecRkESjd26YekUTjWW/kDP2Sw9VryT545RgP0wMU
AWqJaHN/4TCc2a9dCYdId1fwoicwPLbw5HBOuUqFeVhM3zEgfRmFawmSj8DE6BNTcKNGhay0AKOU
udlrkgdGzOvfk3n4NaI6KjRbgTW0dxWUywofMHyc8gyM4lKuYCjM7++w0uCddheJghS1zpas1jIt
uRMeLOP0d2MMuFfr5bxopuY77y9ku0iZktb6yNVNFv5EGvjUrmpiL3huJ9ejhA7OvHhaRyL0bAxQ
9ejO+zhh18A567q9Wj+zp0fMgpc3Xusj7Rpc2dVAylV0qznBS1v1jff6gYavQj633dQrM9FaPWsd
CNOhhBvW4O6SCUzvynglRvZN46I1GE9yup94hKRdmND7Rety88m84rj5UK6oAyLBOnw6Ke4s9zsk
IAHUjVL2syYV0A4IFcN09rAOwpy9tWCeZUr0tPlq5Gr0ywP3a/sx9estbJSAocDtil3G5fOpMhGr
RCOfh58nwB4X4FeR2WN/UOdAbVheJYR20E3VzvjYpTizeasUPBta/b30UkGzjbkCNhw7DwIDhGeh
DVgcwx6HNtGKzZ+9du0bJNyeAjD6c6415dO4rw1qLP1Y9YXaX7LK8DOoeIINjZtn+mUyQ5S5d1DZ
TBXjFi8vI0fOG4alqVzE4AOYmejWevlqlgJh+fo1wB4N5oS1YNOcBvFKPS7vyihNN7HnePrlW20T
3LJ6VgXM8jvvcZHTk+wjPGFZZjennvLSuwTHXPsG0WdfgCdw90X5QXY/K5cYu49If0DPzWr1sso2
OdzUyA6OSyDqdKQcKr9nDsQUsMttdZVdfktPa4JKsZ52QsWYCUBYn6ZaabTLphs4c34X8wkNHYTB
QYhEcTdlw5lxH382JxnmT7iaIGq+ikkaK8ciG7+XpW8vAZwx+iYD4bcsKo/zJ3n99t2c9TBSfcJk
li3BH56WqARrBNQscbTAfhP4HUtpxC4hYuLZ08aIqRx1K0V93rtO/KhDR7oTiZEDxSXqNSaNbd8F
eQarLBlUfgclEZSaZUSCFrdvOgHIWms0oIFuyLs+KceUS7THECHhpzVyo92J1pNc9lQCZ19kLeXr
qpWv5N6PECvMSY7xaztl4ca41zjLaPVAhRd8chs7B5/Z38yBT0HtYIk79A5xnZZnk51k1pNcl32a
Tf/sEANjiUjnavWZVb4z/bzJKEBBAsXoeS9aQ2/X8O6iFHQayNmnlUMgwM04/4qOkkAscCO+qURG
W77zddfBjoNxo1cdwkTPQHKaTcK5fdgnDdSZ6Zq7+DCxrHkkPk0eWuHyvYQ2Ae+Dg7MeSl9u7v42
ZeJaHGaUOKlJUNV25O+sKApm4Pg7pB6kpvn27eA/OVE7Wka5I6nuFit3M4Z0qP5x/ZLEJbrfuLCo
p8Qwwtjqf5TJuT4H79jkaeLr0rjsqrzAQ7FHQ+jwigqqB0rzLITV3pM4ZMfdWLlwq/NI/FeBs0xO
apSkb0xyiPsTYENoZlGPyeNopklEMLVRrrKqK7yt4x0yYOGe5nYLuX2H/6+Sz9vG+VgAoz69lotM
7RjbKbcrdI7rE6zffouOimBBTdUTChqUF2/aASTkiafnQHy7e6Na9/dGFcFJMy2P/n+2Qml98b7C
kOdnDBQMm5bAF6WCul6LzfCSxlcQNFfyvTE0+ZmuXxEkgLlsMCfE9FvldAJN/DzlqmUxMpu1f9cr
SbF6rh3WXmm5pDInMuecp1+56ntwLfpXsgKqpEltmNshffcqTrN/dTOYNfoGAcnfy0+cBQiFlbRr
H9FmIbZJQ98mfI1szD4hFHCd9A1rSca+bxxbpO/67cEQvu6IaBUA0qCxUcE601b80Kg8QyJQjU/l
v4CGLXnsoHhE3Q3nTg5caausw/AE8Gl/Mz6zHUqeib7tMCWYVJodNYBf62Re2ooMFvFwzL630PHZ
W244aJxZxRPp3r6L78dQdMnJG+6zLg8yTjmOr4zuw27RM+HVQYCqGcgEVYfjfLitZ2Ei3M7foJGf
1WrqhkdQSXogLDZ8MwcbeiCBLZukQOMB5VRMpO5jtc5ZFfwcIwCRW+lpLDPPLoojSKDKyNoz0XzS
bMlFKr1+dYQvgiP+t7MNH6qMza3t6eIrnjVR3IVnQV8QCaeT/jt8LjMpFuvvSZ900cuRbrY4DdnY
VGnnVagLQyufEW2AL+jX/0mVC5rjM1VAWxFwX3kXkhvkEPwDP9zZU69Lf4YwfTmmed4WUQ21gM0J
QblgJ3658wRBqnbhh/MAxnkzSymWpcBnPUXIYHZ5AYUx/jVsM0nW/R0mVFXGbx83TvcV4ShmzJwS
p2FO4VqLFbESE9rHWgvHC8QVvdS+VMNLC+TFRfSg9QZ2g2GG2VjL5JyG5/sBgNYaQLjNDQeFgbZZ
da4njODOgiUCxqfgvF3qsT3oOaxybVixJJqCtmBB0nrboiggO900u6Fg2g5OR9FlFNMjUBiH7gzn
tf2omv6w3bz+66fjXWGUj6eYzR/YfNUzGPlR3hUCLXHGLwhuBC6sAcbuD+Y/w8YZQJ9x5cxrOWqT
Jk2wIZWT01xnQHTGRw7iulyLDBaa55G8X6fvwj4licEmyrn4MjQYND+SMoB5UAonuqd1epY9yaj9
FSxFQbZJUfvuCp+tIMmBZJlacTQSSpmFa35scZ2yje/CSwBty3R5DhzbkqQM0n2xAqPmhPf+Zw25
lF5c1U1sYDrfDurJoO7zYi797qE7p4ZxN+0Y6nhxidR5IDy2wyWlfW6aVCvW+nkGQ1cX80NHb9cM
Y0ERtFasuGflM0oGW+CE7MbVHjZk7xovyccEo4oDGrixSZSTdhhWyGIFI48c/4iS45f0rRqHFbeT
vm/r1RUc72c0At2Q2LZbKizGNomFuvWBlTBYaHcXYSxu/l0+fbWlQo4rrQy0kA9bMzfSe1v02wbD
+3UewM3HGD6USWrdyHZFMLs0kn3HKIK8poNqLQL5idG/BIN/NlCnTwAvwDpa5+LQggQ0qRRThkgx
rIsN6L5OHm2CHSgeACovFDHH9oi6P4ioJhC+2TLUVNUjStQynUfXjd6xGvuizfdUInqxnVsDlGLC
JVgBRnaTOsEu4L5CojfsSiCkjo9aoUO48W4ADx7LUHk5o1qq+bhgq0Jnv2GcaqToxOvVPUO0dIbc
kTUutox+Nyp66SqqFoql/sm9QDQatk2Bein1SvZu9bRod3CRGfeTS6kMrgI4TUj5qrRLm78SFEk1
UsfYSMS7fThwQ1gtUycIxHaBLO53fnqOT9bhlNQ2pHQy/RofHO5qJtIHE1gH2bdk4OepIWGKmVoJ
n+ECc7nU+Ni0wVoz1BKSwLiQtDH9H9yqFiSFlwS+J6KjV+A0DBFcyf4hENgqrFIVCMGmEl9QWH1X
KumL6R5K2xeBs6xaQVRHpt4kATWLa9TRyFePodEq1xwzIyH/JfRkDKiQ1my8mPv2OELB8QL1EHYP
qkhYenSoAxxBfcb7fCHs/ysv/Fc9HYmdfJQAU+e6B3iklq0uYDruVybnCPtqkO/dHSwq3RigsOe4
jJIYyWWENqAy2iDwapnw5NJmv2qAFfgoo4EU+IsWtIui2wf5dwePoGdlpf5dtrA4z8/J27b7JUZs
w5oxRIpUFKxF/ozq0fMKls8MV4VN1Zu7dhk7A92h2UVS0MYOId4tXThVcWj+h0NyMAoGDVEUzDxX
9khNo0P7CSYJtR0D33Hcg7ZB176Od8ty8gjfZk5MrcfoXYjf1bWCnWrrCvrVDm46e8gNRCVz/n0R
vJrZFyOSycKWPKEiC+XZYCOfYTgkbbG5Ms92ylBgUrH2okMdvPXWsEFgzUCQ5IIZjhRvMktbYqUd
kAahonEKvPzsD/uKfJsfkz/fQ+AGCPkaYdqlT0YsLxpjfXNqgyw6B09Dslb9T24vo4U7t/b7qsuD
ogrLzudkl+LIGaRxHkoTN2+/06gUPJlO+giiM5e+62AvO10c8n4UCLjmAjkpQ6hVSpX+aAgkS8qS
gQWBbKbHxKfTrEQrERNnaAOckdtyWRQS06F0AzTbi7mO1pGqjiwTgcFgFJMPL1upc6oC7juF4nHU
HvA+ANqZXJjMmiKev/lS34XhMEXbhvVXurRJW3moM4Eew0a3kuhrGoKsAryHUgv2IqKiopHjSvY7
oQiyslVVsDekp89LtnrVUbPxen2pEwPoiabSTOa/xb31yD6/l4NL5DCebBrRzkXd5iVbaoZthj4p
MfbVAccvCnlDjItvnIe2HG6Cfsaqhee46XVaiOJoOijKX9B7OggSZeVcDKAh6EQchmg1ZluWWEMG
NmtEX4MM3VSlSg/rT3pgpR4i2Zxq3SDg27vXMz6jserKtO+yPVhuh6c6roW4L9NUDATtji1IyD+A
S6rgD3GWS6qQZP5Xn5tU9hvBB8JmB60C7TTh7sXVicbfKxA5IaqV97QEb/RFrzhzsrwX3oSYzTme
qCfDrKRgrQo/F2J0dxVzc7NTEhcy2GLJ+Y63h9YuZU+Wby3nxpAurfCl7mzBssOhUC8pVyGK2ClZ
+DI5CsYryh/bX6MJQEKJE04Eg5egoNLH7Bjo9IjN1yVh3b1rhmgmUMbkzbVWP3pazajSd+w8a7ZB
fuyiCHiYGtwAwfeO9CIOtykv4rG1zvScy5NrE5beHg9iun5tt6OKEvLYjrwMTqAe1YhwfyUVqokC
k5u32IelJZspXF/DdUW+MtAin03c1rbEc1wkDXF9dGwrRpO6P6MbJPfmP5q1+Ijk4+PXbzxffQbZ
hN4VET+ue+HthrpqtTgMaUAQtzKPXPC70U1gCWnUHCrGyY9kVv/ymvBGUogJ5lHyk6U/kZYd1ixc
jpKXeHyIns6x6tB5pVx+g9lgfHvKrR7I8gVwjLzoWMXSE6XA4VnBQjXpQOuEg85EbN0OmlyIp03k
rzGUSCT/V7ntp5iMdeoXeyWui455RtrjzXm6GaCQT6mT0VGF5HQFzXxty4rM4OiIpvVZfy2DP6kx
Hr5J9OFutE7XlB6IR07JKi71fnr9bs8lcIqTwDt5AUdDYH/4uQFAa/2y/ht47pzGYo7ED1yIhkar
inuI+jtq6/iaegAjHgu2aOqaDcPZW/GW/Ziz6kPAaIekgi9gMZNjTazntGXokQFZJS3ku2vD08pR
FcyNQSN9Dy2matORMjAgH9jGPAloR9XXn3WgOrG6BdS6ZsyfLm9n7/4YxbpZ8AvCfowVx1n91y9E
ftlEebAzA/pThasalHeeuybMpoZuku7zuFNqyNExO3QCKKyLcmEsjAnSDT0WqZGoM/Qa2Ses1J9R
RgJJsUEAfsgo+L8YSd3uuq9Qm/FgLv4gmulUdZik67WalknV0tRIUV8QLLVaTxQtnGD5RSHhEveS
OFI9EZs1sZEoB03rYM1Sjw4lM+0RL0ZfyyVvaTg7S28Im2PgV3fhjeQSsWzoMuWtJt856Qg6pEo6
ab9+FtLLrOQT5lA0nyNIeU5tscWzm0UZ9GAlY0CIju+D9K5nWlsbmtV1IkUs5N6w3TonIdS999VF
qalypDtpe/fp/f+OFetFyggR2wThvFm+9MzcGwZy4p7mHzDudNR9taNaFn8zPQZsQ0b3FwdSSsPp
fdpyWom/O9nVGfg+qMMB49dHYRHhOn/bmYAUPnEDCuuoGYEZAyF3XAzS/xDM9sWRS6sMsyNCjef4
q4QKPzZthXYgel4vEFomj2R+YhkYH3hUYdUX4HBtE9tUeUcjdcyKe+9YArgoMFpya+mTj+fOWkcb
FmJPAryUr+yPwdAwmtvuXUFBsUEPB2+yLe0inIJ963cJCAbMW2Kr4tokZEGSiprsugR2LtYHkH1X
9j3oayeAzepmsdVkVDm4qogwQ7qOf3SUkTmkaka09cFWWRlwpQ55jJKmsLTEOQV/VV1litBGe7ZR
4qtVv3RB4RqnVV/itqDoeP3i3Oiu4NjR3dCjOD7I7mE3itvm1h10af3NFMBVBP6zmU140+WwFqoU
rd34E5H1LGHGcZWaUMbsRtXmBVXFxPCrrvrG2XmYu2GpfABl97ZYDqo2jjKEkIdcUaRwwjPcEp8S
jFVzmGgEDfUBPDzxqpv54C53lkWT7Oe+PIEQDgv7imfApnxZ0mEdTGLgF68YOfc2bed2AzVGNQo5
S7bhGdg9d9GCJJncWBNp5iBqyBLRMez7AKEuYJAKAOhBNEXbLsm6Ei1AiBC1YL90qzDnJAt9OJYz
RHmFbiQKbcPJ0Qo7slKanqQdVg3Qz+NgblJpj8MhkBLEy2nzmyltsheA+r/D6OacMIIT6Axsugdi
CsjScw+GnRKLvuOOuB8pyoKXXFfbpdpka4u9X1wvFjnR2ctc+RYOwkd26v9yHb7TYS/bUi6zAc8G
l0xHlqSAHt91PQK+Nolp662rgPnmkx/td+2i7gv26zBdRj+cu+5VfXNoSDE/ZPABlVsYy118YRpv
khvHKhuPLQruIK3uY7VJrZ8IoejvVdAIZg09D/4laWIoVKIL/iodCcFWQeb2hiSqXVhVOVe6p5cb
1CfLHNf9nJhv/82ZIucpsfK7TQrHyv2ccRufNgNmBuUSgIW6NyS0FWnbUgIhy3FdiNklpJpUB2DO
OcRJqHwBwnq/nCaXeY7BYO5f1s1QwdpTyOCadn4SXM6+NGFmuKrxA97FwjIxyAG+XY0NKoKu1VqI
JHfG18vH4inA4Qd0qsabbRU4lJ4g9IgvqVyIArBkJhnn5OliId1qbAttkVdBaPeP3u5Jiwqy6Sff
oksqVr4WvQOw0OZfnQBSJouhn29eBzp4nvDv0Ws18IguRAsiSuE0QiGjRK30irGfp3mWgZEbAtIg
qY0bzthZueLzhxXBanCAlxrVH+UKckQXoOAHXSPdB9GrixI988HbQ35WqgNuROdJiRcgA+wKVaVu
5JFJy+XjNqVj5IrUqIscKIbeNXIdU+YzlOOUoTLVe1/6Wcq0eQvk9WDGuYRmd3kkdcgp4WbaP2Rq
n96OrgUelBDfr6nWt3rUFXwk572LZVLRB7ZgmmuR8Xh8XiVkULMGQIur7IA4dg9lul2LpWZRQHeH
ND0KfjUHjousOMa/nPL1W6KEnmVxcCdZvzsGrA8XckOkiSVIcYn76ros3M07iRohZu6VUbR5LOyM
Hz8K5FT0O26UUemT3wyrr9SCbHd7WKi6a90wiqqTpYNAdbzhwCaaNygBqx7+zDdpGfpr3huxmSjE
7wzlopB39KeMl0ODcqyKsLpAG2I8U50XbLcXbDBIZ3dKWWQjz9ZSPVQdzqTWbIraQ3WpSM8BrZlM
taqiIyy9qOx7ILJ1l8jvaows7LIEIUnAf8U1c+Fjc5VbLlvyEb/9lJ2BKBMLL2ldjAYX5efoGLDm
0i9qCOExk2vpilz9zet7KapHjYlfxof+g7GwRSso8vvviouQZBfS3msi2KbFCDAkXYWiJc7nuAEc
BV5qvRW7WTbfOC7ObtYcS+m69POklAQ992nZqSnranCvODzLqHqsCPOEJNcBoHaPkTXbJSD4JCkI
+mS/QbVNfsaGWJxKzJqK8lnwPag0uMfUOTw3tj2bf9h3TkPnzuVJykfUcI/RMcANMeR2dBvswG7B
uH35jl59WPnq4Q+nl+YKPisQQExw+Zv08OWjaZvuRbZdwj0ddE4+ZxyUNl9FXfNeXfRKwwf6gsbH
47XiIk+0AFDDAGUiDf6gBjdql6i1LdN6wRqgU96kNdCXOiKROm4z2btkzspfMy13DxzbxDUa1qKP
pDxKzq6RTYZGxG1w1l3OPFn/Bxr5/KdVq6+zYa9J3DAzib3vNwZIAmv1R6bJIX9Ea7ijafk02na6
KrattvTmmbjHt9f44e+O1HoV+1w8YxmwKl8OkKcknO9Z0qbzFxn2flOH4x+3H5RdZ0yDsQSwPl+y
OTJ10qQcs6X2L0EPXs2KdrM69RYf+LV06JsHHBmVttoMyLaDkj5d10ta8c/aaA3dUQ24ypT4OMXp
AVGxLHcNLPK3czsQxkUeVb5yeG4hPik/1R0mEa07OMMTjQfhXp1b8p+3YGGUPr3nwAfJHhHBXKfS
DXmsOpAAVVbD318g74lmMlNQpM6U7N0ZxN55OtxYiHOSZ6l1rWq6Ggh9sr3NJuVNbBRAwvGI58Of
X5W01s4in8h1dAPMSE+vx8MVs1VnnsX+DdACw8z6bpj+V1DDQAoXM/fwU7/fAuoHdiHRoe+QFbq/
nD3svONTPti8TCjS02yznz0aG5tUtMxJmRZDUkDXGOcbWR+S2QgNOAmrophdFcc6FVtuSw+ADrDV
1okHIZ5bMxmgeRG1tnff3spToY5qo563W9x0lX4Rr5lqVuE9JqqHRZ1tvp5JVe60pbtZFoCxYCQH
FM9ODqrF4p3IcqTOvHg1NJAk4V65jjjsJwXrwfc/Oo9UFoFJlGCooQHO0VG4pM3rE8rNAiyDwxfm
J1zBbYjCMaQC/sjNbJeKJFx6hJZkJ56Q6y+UeEBgPeh5fz9MDkzfA6V0m099Ww0M/oNnSv3AOhsp
xqKMUhP3e0vEkavrgfKM2sizt9326079Vc3CDn+YBiQ71IpfWgkwYJsgJtXX7/SFFXddy4MlrxVN
n105MjMMf+gP7xR2lYNcRE7WQ5VTh3gQiqVJX5wIF+65UNfOMJe5fDJIpc0nOVa/mVOiIm1D4Ail
A5eX8ydKL3yQRvRTCNCL5Ip7LYX6lVsO4V8er/YCPgsROdSZqVoZ9GaRGJIm1kSA7nxpIPsyin1r
/36VKT3+GAAuA++5xwCI2GGgbhn9pOzcK46pAos3pDROHUm7Hxvnp3dCmgCsh18UxRETqDN+o9FZ
+EBUrK8OT0DRZ4zu3eg9gq7Gi3ZCr6o24bpAu0I3cXrXtp5A4V44rtySEvm3gDp4XBLcKGImtq8a
HLZ454EEYzJYaj4NgRdjgEleBkD2TF//TxFRazjUjtcViPjgXNH99bZB6ZbHQvYU80BI/Ks9fBy5
VBzxbe0gQJE/mSr3CDkWK4cV9SEbNA3a0qQJptEJ96wMJNzKThd3NrXiR0KT2KVVIXmTQt1SUA7r
1v3/bz1yCfsA2m951Hs56y88Ivml4aQN8NeAqc5enL7aWnqanvyw2YpknkmX2g+4dxneVCSDn4Ig
43YsmDt4MSvf0QBA1C6ohQ46VIzJQEqBBH9dTjpVUFxZnhZKe/QMLnxoVaNsXWosCLS7zdp82cIS
QqD/+oip5BLWSDKLntRw4lKBQ36VgI5g9vPmBcJCYVr6kBs5TLwHtIuulhI1Nvfx2lmrzez/UaSc
J1SNfpMKwFO5D/FJNR/PEPy1G7ePS34igB9tLuiTOl0ksyBt71ftaAhtjYLDAecjjBGhHslDfG6J
q2VLKlqr/gVFw5lAWXbJhekcGr2AUm9O5eqJEAR890LEdDOoPFGKeYDZtKZ2WsmFsPFliawd0P24
wdVyM+wp9TqdXkDnFXWyX4uAUjVQGT2nESZ8CQ7EiiPNE6l8jTxC7p2rKElsgGLBuagMshVRdIJp
jFZzcQaK8/bb5DxNQUyeqFRQLDtWTwSJf2szr6IW9wfxxN9It9EHlxQarnohCt6zq7D/Enz6gGjP
niW2fUfAQ9WTKVsYHcgi4ngnOARKELSkdhqp845QuO7oZGRIsCxG5a4JxlEof53bIS1rbuJQKnNw
108zzGxTMf5elwk7KoLdBwHszPu+muUx/yVnbjkdqIXuTTM9TopD8znSucDiDG9/hGGSmeqMH4c5
5DBfGAgqDt+rYFf7RvvZ8uS/HhX3tcX5yZXxHNtyp6+OonjEbVdEcF7TSl4NcgSuwqu66Oj7NhD2
2BBc2HehmZmdFSTB0b+wEuwsxv/cS/ISbhvbB+gtQH6dqffz1wfKISzImBE0yaOlPMJOLZAvnVFN
CWZmTa3DNqgZWO33L+kP11oQe4ps/jrtr9gKuzlr3uvtp3dwNawZfNqV693q0KmWt+F0NYqEd7gR
pCKmViQmEDUwtsB2wYMQR+rPQk0WcEKRjNWvwP6u6sc07Nx+xRwFPZ+UJI16WkcwO6eE3mhse5KI
VX8hO9Tmzc2Ublk2lJrTOzBmfKyWtKkDmUKrluu8hLW97V1hTDJkrNOv5KGHfV7Gyz3dbOMNB/Gr
NB9BKojrWMpO8VvwB+zxghKpT52cEkYOKN8c+CE2rB/l/mdJyLllZ6a9Ls4I3tmjm7/G3PmfY+2B
Vqnxa7z2zyF9rCB0KENomueVuQ/1fBv0/amSyWVkxGf3Ym60fKc+/h8nnKSSUXwLyxHZLCXrunAz
iLDHNnAHrh5mVZuGazdPFQ7Ai6qHI8eh/bAFfbaGF+CUXsdpK4N/HQk6qT27c2ImYCWWB3qUO/Ln
Kupv8fIkdW1KG0SdXxUU+osyAnoMwFlfRCEKFWcYPlap/NJVNzrDBNN7rL58Kqh69LtumOwBqJ9h
D10SOMhCa7MdnJU4Gimi3Xh79xju9yjsudrV8EmLS08DmRQhmz3wM+4zYSksW17VZYlKjbITAU/X
xuFKyHanNDWkSmgFR+m5YffAAQoIPHrQBINfBfEHDaHRZh+NrZKDmiIeM2aBsiT/aYyqQ3hpW5eL
crrhnjCEJDt9EVHrgxIayd8YXBeM0rIymDzuyWCtk8oEIQr6+FM/ouEmFqUU4jF1gXGiISSGvhBW
cFZDBGylb3Ff9KvBCEPCzCHKW3FkmopvgPAGcpiuVa486bCDJ0vsjTu6TY2YwUnK7gbJT0bQFhlD
jhAl346MYs+vwz1rxFuUMz3xg5du04zm39a3o9MPV8a5l54z04flNvDB8YNF7CMOH1KYgxWEa+Cp
Dgq+l4ZzujxVWnv2jMpipexBv3bdiWwfMQsPVXMa1xIoif/PP17wLAW40JC0rcUZazM1M+eJfzpK
eLxYAzCXgiS0MOokaVfiYm6/JAZY6RUvckBZNgyZaQaFRSvQNRgb+rg39pW+2LpfL0Fp/nn1SPX0
ix1D4QkQBHRpEFync1FLTI4U+dP0noYHGuhe9oDwH+scK60de0OJyJmwvRH4Ac9+p84ukizmgt4J
PLWXdRPBhsO7N6q0Tr9RrHOB9NcWeUI2z990yNWZ3mHmEiv+Z3vQx+7fIbMfE/EiuFR7FOwWbSus
2W0xp+wecexVyIIY3ding8ASD4FwSDcxDrP6um/rlZg5ctx+KPBBuEN4iNLV7y7OvTPiOl4jVL+j
5MgbBQX2AY9m3njNI5XgWik1lOX1xlHFRcxoxqHTHpkpkOQ8ya0hKbF7wb7p8BC8DIxjns7yr+6z
CSdIqG40ZIBXtJjY4nzX9PitB+AsQM9/QuPTBaGNGEF1wju3GrtL6Rpynywy7ekZt5cgddrf8XWg
6+1m0BLwLhTcPR2REi3iupj6mLHlSwhaVMms+IbIm4qA9Ri8175W77Mo7ZbbNJBoHjE/PByovTpK
mQYVQJQpiHLbjL9cjDuIjUU4R770XZEyVnE8RPWCHyMkIvZEV6SRDoo8aZMambDN7Hms01KN2/mQ
hiKKvh2bPew4nWFm8pHSjqNvIh72FyGwIxBEgORVGP/buEjUIbsSiRCUDJtrD5IPr4F2i3pTrFLb
cqjQFZp4tTdmy6aMSX7ohneq+2pm8Bdl3rWA49cZOQiuErKH1Ap525UK9lW98/MPR1XNJ2/le3Sr
Cgpbe4KqD8jLdq8xXR5N95FKvsnZbyaZdELB1Qik+1ugfCzHy3MM2XM89QVMTAsfouv8jn0NXnch
TZEq/dygc4Dca01DHAWV9tbiyosCrj78dLafMx8PZMwMxXBhzfZH7FyAbHK26MtH+396ji8ECeAX
z3M3PIrqYhmhUQZ0M+Ci4SNQH8JKywRXCO+YzUtRga9cM644QXsSIVMF7zDma+9eeSjvsQIyEWYN
8JmzX6jPvf23/UofN+fSETQeJuAFrTvU+a/1dV4tSEFU6kB1D1oFUMr/A9/b6Wi7uFAVLshwwHy7
fdUb0pgDgDeD0vhrL1q+TuI4AiALlQZ+uD3gNmVCf1czJ9YOEnGWSQi0ZUlhs/16JG/j3QxqTQov
pCcev6xSokN3baZqdbqFsvKsgwdRXHvn4VRFrVcBywJAiah61BGEA+eRshlPxkKFpyNoQmRXRfsL
o4PbyKwgeIJ/9slapPZxcREZr4o8GqVgkDekVYzsE9OwX6MI5G4DUqcQpi/nM39q/K8Uq04MycO+
xaG/62TAeQNr/43lMVJbfhZ1NJ4cmRYdro52KIUg6OGfL+Thb7Vv7zso+muS24PkmDFUoTqayYNR
hM+cPL2yUume+R1XMEziTP/TIAYdZ60JbX6u06uGe2lLS+MP50AkaIO1eC2FcxmZpGcYap3XFQaD
hnvlP5xdVaPN7Si5TwIbhu66SB0hFoeEMMRzAx5BbGhaWCRThzb4D14cyoBQwNHgghvecq/UBTSK
ABP73Pt4DULze/UWoEqYNpmJ9qAlTbaol5C0IIUbX11O74gaHAWMU6JIaurLIMY1i40+ub22Yks+
XXbjzIcPRt9eSaq8+vFETh4+/1vxor14y8rzIc4ZbYdCxeBMmr/JSjeLmfo1vVuq+prVsNaB/bUI
/c1JGz9yewS/9ZWUI/l3t6BaQlSfTNfGV8uTKJMr4mKGb3YLxKnLh17dyw9vO/V44TEsFTPdXfC7
bMcFjm/8sD4cQ9eitge9xjGRqVN4yDtwMMAUEPEMERIxbWQPxJIdrUZgNBWrYPAtijgFN/BPpwA+
Dd1XwoCyslraqN8BV4/kyI0wsRKpu8ghG0dXJNSm/AnAPXq3jplNYGb5J2FLexI0YmctweVNMdRS
tR/CtXRUcCrTjwVA6j+h8zT+SIINVIJNYAKoVzUPSd1/vYmVey5i/7ktWtLBjd3iGxNcVVKk5Ib8
ycnh6IW7D4SoPfyePSnTCGmS4PP37i4NXSdBxxahlBVr5xV9yMkueS8WAdY5kG/6M36DAL2arDhD
VewsjMHaJTOQWu6jILmaqQOAM+bxfB+yTta3pSFB2RiKo0ONy54XO+QK2mlkdbfwnDWBR6peBcKH
J9nrywjN6oaSWCTvTikw8Ju33uMxozygxkOADutFgRcMDnmPtbJaO1u0e2ArSBeSqxKkae/KkKFA
7J9pdLXDewvUKHkJgAVx4BF+eij9JPrNFtq3dugkeYSYR1tsx1BHLxqyUC+yR1cpfqKXzp9Ar4Hc
kYXX2TzPocUA5B2XkOVPfzMs/6d0bV+BtnjwCb32h0bY/FOKJQ/8JZl1emis7F8dJcKEdqy9sX0a
fNOk2Gd1rddMDCh/JjZJ4CNrn9oxpR76K7sWAsYw4ojeT1Kp1lRAAlYz8oIITb8zQoIRfOkaaEkY
AHAItw1JyBv5pG/0sMXVJVVvaC+ZMgMtQPAzHuQlza+PvQlYoLA1feDFzwmZLBjqrSF7et0YFsQu
za2oVlCFoCeMSTbX3DPoW2qihyKvFABrlPDB1alPB4XqWrANV3zfhHHOVqv5PWEKpDPLoNFJnyDh
8e//6WB/LMZzTsEKGLgKzs/tFedpilUEJ4a0g0clQCjaNf9QPJg24Aag4L7nWM7GExR2Ezu0xuAH
eRewlSKbKlu2kXz9Rv+y19VYVuGAmnpBu0Ux0rqlsXc2EonBb3CjZvXK3F/7+Tt3GkyBuBIGFArj
GvVBpmF1WLomcsfqbtePka+oRFi27uUaKONh7mxgCwp5mw2B6PjsdKAYPjaAuyc6FdxlP2pBXqDN
BKDp50UA9Z3CkmTsj67Sa3zxIEeun+UQp3NVHXyOaP6XNWHIPRh7sOy3Ess4y1eDTUY4HDux2gf+
p0gWEkJ95EEcySLpJQCXWWhbyaxlQ6clbqmZDKc9EYy2E4bnXofIZoRJ2Ak+ZXjJDcZLiEwhz0/P
xS5jrE/8efZkUvcbXXD7GQWeYlM7bivE7h9+z/VEgfziZT3AIFcPiPL2PYjG64i68qn92WT0qXY2
C4zoBI8kQEpv8hEzgsVBibhdhL5FSesJpCYvnJNcP9JuKM9BZ/1FcQfIY2kfSk3RbJlw9msoDGqL
nEGzM5P0TXJag1G8xUB/JuSLl3XFi89o3jq6dP/hfoIPeiQHVrvsw2ZZFqmtatqoNu4A172dL0Aa
DLzIsBBybaPmCa/+CVIaa/Fe2c/Isn+onpLgDD33iXD/5AqgluXJqGNYFGASofS5CupcOBq2+2Rv
IBfnzLiDSSy/3m+zMH0D1dE7mlcI7ZZHcGDsWU8uzcA6NU/FI551bPUoP+NxmqmjOkctMogpk19+
2zdd3HzfIG6iDusblUh/UMYXbdWHymmRb9o3nJmGtGOjguitCAAYigb3dwYORpF6nXoS4swyzm+X
JiVbjQA9DhIrdg8cY0o9PTrLVLkqHcgdV93Jx3XCnkUVZUN/CrM2ialb+qX15SsT110jYvc0AMhZ
Noh85mpCnCUbAHVJ2FITRl0lYw3meO7MIw5xg3NX2seS6pKSXaOB2V+tsPRy9vNAguEfXz1gxBeo
O/jYfr55r4VGwX+lJlSTM8z4ur0xuVSSgmaYgQNoc5NgAkrYsSRGh7CKfltAICaoO7/fSg3sHlJK
Tr/VkgRDYPCwMSsM3dLHF6E8WytlhUELdMi3+VnO5HJsu6ZuLt3JRCjyvjawcD1gNvok3++CNKH3
W2hmIF4JcUupxObquC31kLkovIdIHrfMp1CfdFh7jqmy60264vX7y/Z/meozIO09gXY0f+GDSbSX
WYMFuyyGX7b20qjB4lm4fbfur+wXVCbF2JTOzQmrwAlIUCh1sOVkko/JFob8yCu8I2MhUiWVO8pL
MmiNjydlYhlgAccNHOaiORZRDoRmDb7lhIW1T/wz/qdb7OBasM69LGubvlLMVi/Gu+y9FDl/xm0z
1wu3HwdwDX5zTq1LU7ww/vT9Mg66UAWDfdCYeK23+qomjXMoUkgPtf26mPv8JSxGVA6MGilWCp84
vb967J5+oC8CWLBHw8dW7SM8cxnRqShPfNqQBKBpX4pz0WmOaeTMrSzM4mhV0Q4H77nARjlNfPfl
AeQvVvVS6kRl3h4+ARZX92CXiEaz1Eo6hM9EJfQ9FDtV1VdVPNbiLJouzMxNQpqtPEVYRbNDb9Da
Ojw8m5bTJyp3wavhFiKndIA4oBwWRj8OoVQxr92I+zBDFhaxsUEOUTsNNt44iKRmrYJeumB0tyU6
Vok87jnpyYzHB9sWs1kxL8GyBZhZsl5rcokztighxHhJuc3wnfu89aak7cBrum8XczLZ6jgQWpqh
PIFIV1K8RiWqD36WF7J5aAa+zz6OHatNaWXHsFGPoiSmSZTPWnvpcEaLQMJqCOR0MGQl2Ci/pdxk
U8R5LmwiMU8w7wAZ4r+gRu82YB7jWE62D9bjxcYdkemIdAWtIVY6uZ6S2qrFOOmjWLuQzHZ4g14M
ojxHgzehU95PK0CTfOrXGTlIdegtkbEZhcW5cZEFclH5NPV5AI8zhXaNlD5Q4zLv2d1YsK9YqeOe
cV++8XqfGjCk0w3zbpQpDmvJ9Hd2mhOP5uROmGdS/8eig+s7hp/yGiYeC9ShC4aBuUWIBOCwTopg
HD3guB0AcND0SrgyHVpVGBovjEHxZCSzLYkt2x9Wu90Sypqv/UylF+VYFp6rzOAtZ6TCFgQy/81F
+OpnKy9QCXvMLGv9QzZitX49oU6kW9RBBipse+B6brk3cMp4j0BMutUwkfsnYMv52czhmS23KeGu
aoO7cRmAxNZ6sWBuI6xM/jQeVdNJYBQSleZLWZb4cMqd+OZnxs68qnosH8kXpWZHo2v5LIgvEo1N
KFyeV47IybK92EVihNQApttJg0wXlxRu9r/pzsqt1NzYyiDE2wBspRJmbIedqPId5puTPWpsrrFA
eN+OqcnqgkyoeymCSWrBmnJbFETNgsJ4y6KTea2QxKr30NiINVFaGTHXNZKC8M2UrbPTlhS5lahd
uA32q4Q7pYU7/u/AqT9y1aGQD5ylrNlQULtc6EVfGyCnfAOUu8RWazu9hwVaYqjo2yMEmtKLvJUw
ZVkw5EQvRz96X/55cPb6vR+eSOD/dUCP1gwovfxpfrHHnWBgU9Cn1TCYCJnOoRqlVfUAGMkODsxy
3YnDzUH0IxRUy4GDFCh52MahSrh1TJ8EhmrA0ltaaHMl/gJHD7AKFxxsdHDV9kcKSdhUOgGaDN3i
tdGbqccWkle5TGugJR9S1EIbYNvGFARaCMEjNwpmck+ihJ3El5mU03D7YeZK7bMx3SYRc8vz/bwO
AzRjgJb6SLMDTyNN7UXmg83hqeQDgOFUjKy07zlorIo6/1KMne2hkuti3LF/V3IqcrwpI3iywB0T
h+WN7ZyodR/nG+FqTnlozfP+NWmnG0zr/ukHhW0EviBVLJsrey1SIpcEyvN6wuLyyQAOiNFEZhk6
okXgzn3hUIobsI/lYWjQKywut+nHMeJbUNoUHw3ADgi920L/g6Z+pDZYI7Au3mlTde7NHMIz9k92
8A+jHsPOFRqCVVenpzIGmEK6zosZ/PyR4F3O0ETKKdmcBGWkGmTcQ9VXMKnoFdeUIGGNnpN5NkxZ
46V/pi0KgwR1JhLIqaUmg2Ml423G+1Mg+Z4HOxs76xH0g6tAbpsCiaSSod/J8HRTxDnarJ3mHV3D
DteBJdIFDlhxvYX7YyI7rQx2ihJ7AaacHLCp9pDhzMemu6stRrHQdilz3D4kckGjw79l6iVSs8SB
EhU3ktWXXtBfFYCIvG+KsPS4Z8Hl3rZa2mjTIHygXLRjO1TFlor4mver26bQ1YqvKxY2+wZrOYmi
TK7dLgX3tqqU13Ec+KvcrU49jlq+IMqy44mAbgxRCqeeqfKjZYy8zwQHWUNwhnqduWxB3+4P4ke4
L/67weVAwUluNDow1aPov/XWR7LO6bP64C0wXtdYng+4WUoNMi06yONrAKcJgRLZAsfu4CYgrJRj
2LzJagborJ6L41rajVxXffu67fDg/T89W206qJupGya4OwRCmtBf/ZtrDNV+sJ7VV5VZBQLpQKI/
GXBRvtOIBtMaix3tN4cIaMjXov6ad8UxXNA5GUA2Wi6AA8xaNjsluKSBOjSyHGNocmZR+5WyVJ3d
qwfsSL0vnRZx1nf4jBLW8pS9xJl5SL2PnM2Tpq9AfUUGqjgxrpyu30cfC6di50jr2bNhlJKIaMJ+
P6IZGdPmteS+5r5HNkeCklA/1TJmXuvByoCAg7rdwysc1guU8Z4YV93McotE/doWYOacwaDw3/uN
A1R/o9jr+xqxqyJ9NLnh0rC03bbB/ThXhs1wiGS8gxh6bYU7vJyIbsrxr9RqAuzyL2bcEb9CHhCV
aGXuUTLCR5p0o16DBmrekNORJAZdp/ARTewobm+LfcWpwnOfXkvBRiMdp5AjrU6H1tPCHSW7x5Fj
B90B1mDhR7DY24rCycVMmh+T9linpNrdBjGc8jQcVpcTH5lgFfFwV1jJ0pHE2Q2fX1tkYUgmBgBy
XtlVD1GU98IV8ocOYUSrprkl2yULa5hHPdtZc8t/wfG8wZRHdwRLSeq4J1Sml7+WOx7bj0BP1slu
RCGZUhXYsz046ZOwHqcf1HdktCgnThbA1bom4V/vdee5in4z1uexbHg0cS/0cTGAfWdu2l+1ZbYL
mkFzzkT3sWDI9ZmSjbrPRdWzk2rB8EdYKyx/60ju/42dExmqv5jpClbdJi2VaFSjlnWfBduOm5wy
1SvRpsEKyRy6eKp6e8BTVPB5oW5hKc+tAgWCCqtVqOGLxQRwhoTmGQuS0XH83nMfcx/Lue155Tsg
SK18eIG5bTVMl8c+jljv68oW/bY8jvhdY+K9EltRFUQPj8pWL1j1y+tpnryzMdyQSc52cT30zocj
TD15a6KMlPC6aS59UGjP2c7LSgkwJlw3W08KXLUq6SRNjbPyWv1bnVPg2Z0lzWrehozwubw55/50
+DQwdfo3uYyBzUiYotjbYMpGSqrngAXaSJ/HVIZocwmhq5HobBs2e3LPjWhg0DOurQax1eyo/WV/
21FG3q+f6mU5+y268w8nPJSRAGjUkaZcNZD+RQ8JQyqITQOhEF9EzvrEjAjJ0yTvDta3YdD6Hdvd
LmYhpH9i54AcEWdjQe5YjOXb3UUS4nAqTULjj/yc9qcwG3pyBWcmF4ZYE8bPc1Sdu6o0TSxflMs/
zBENrvIVpxBPge+dFctB9BjEFzHOqf66fMtHiCUK5wM7hzLiCc0d0W14xXuUT1njaKTgrDByFcEU
qdRx5pQPRUc2eOTyw4nF1sHqqnWaZ3CcgfQxRbn77dt77hiv5/IRBXowz1R5Ao/QueiRwTCyMM/6
oRayTquR5Sk0tF84j2htxnx7QULPvXF+uCLUNeXlGH9+mssyUi8tTG7cm2Bl4uQctc7xGLOTrLSg
bZWec1FuZm2rxcsZsmjQxKb30tqL3IIzZRQaM4/KTJbxI/cG7bUXalRuhlmNjmUlqQoudiIVLYyz
foeHDvBwG0f1rhEL69JgfxoDipinoyDsH3rtcG0fSWs6F/IE8iBNzeXL1XJ3XfaZ2wt0zu6BhzZg
WCBlCgr5dEnpv0JyNGDBMnJHJ2zx+QOdEBNBEf7JMQLqGrG0mt9SSAkBdby3US7l4GUuoIa4xjUR
Dist137D3v0WS/2vVbu4iNSbjUxstPVYWXsTWl1qmXV90aNQzCeuomQdlBs8jRr65QlY+eHSuRPc
zaXMQwxEN4Yojr4gguVrkYFtYvpKuu2iAkdYI/jDuxoZL2/wb8Yz3PHeXahivgPRTStVS1U4a87A
lmHKxi7JLyDmD++kBawegUhAULnp6XdSX740j0E4rQcbWaZNGKyVDLMxo4IT53tmWbmjSNYMa+lx
/D6hAQxT6UYh1ziCONYOJQIATNiOvOnhNG4zczVcf8KglcVEP9sB7im1NNjClfos1jfHwj1pUWDM
khxLRdr9eYiztFY3aBKeP3sX21cA7xPE9WoL8GHcw0AcMf8FE5KnEEgXHhou1V3CrAJwEjteGXjO
vlCLYIC77shiKK0IdENxgUgy+WRx2NuxAw4vogBifvTFveSt/P/XITNa68Ktst4jso+Dxalp7cCu
PMv8SxRsMhmXtek7h1p4YoN7wSdteP1i6CshPUPRE0Nji+JFjSVEmAb7fFnpkBbNMnyun41zVhsw
iXFJPpzgwQwr6jE+VbSySJ9rZmkuc9wm486lmt0LIrFt02Dal9Kfa7vZg0Hvi1iyjDz1s3PWH8m9
nFfuSyj5F3jAIO6oTiug4uvEsmzGqNgeGcSmZ+LggSo6OMxSpT0iMYYMiBrOFneTe6Y48S9ePKrR
Buciyi5aSfJbMcDHwtaVmiaMMIQl7OLAL2/UNLZifR7FPjbt941WCM+D+ZFu66HNBfY9s8qt7c0y
OdPdhF16dHRyuU32EQPp+hCjmjWHLU5Kluqvl+pvX+3zj6Kbm4f+Ay6Kw5ypsANUdyT0nPa2ijF9
5llPqTLlzh+9+nNZpjVHizANK1r8jwEQNQj6xuN0WwRIpllbxpChjY6x+hvcF0xHv3JGDJ3FEYQg
94mlTfDnq69rAqj53fdyHtaFL0aT2mxXaYsYhWLTPOsJxJYP63FVIgXDO3LaRZyTptWeY+ej8pKl
HJcTiAATmevtFzx5ySofOcXHrMM8akdHOj7KU3PMoVJZQPVO/U9MHBXyJCe7oNvX7NIAx+D06V4z
VExyHo7tiloyQBs7Dy6g/mPL+bVS+MzEfZB8AX3w2MiSERyVFPCSSyDv6/O/VMgQcHH7dHJ8no1q
mH8RyYoJKfwWM9CZg7bIqBKLo0jdzHWVrcWcbr9Jnt4uHgeOD5hrpqiGUo5fFK7WuqEOD2v39Way
tKcXoU6DVazWpnHZ9LpjqkV7ZMnJdQB0SqLIUrXhUK0dFBT2eajEc0uZfbpPsfDaouAv64tCOXnI
4Rj8si6ozJhIHzo0sxxgSTag5mmdjrHiCBaABDPUJDo7geQYFYJ3+Q1ukE0kUUCUJIFgXfXlN+uw
zI7pGe2dfT4100SesmrpQOCFzT1vsJfCUuWRIJSKPcMHKJoDa9onUv24jI5QbQtCJBiP7xmsfa8h
SoTtVZGzWQqa5CHZe6pL8dMwI6MDFTI362kvmVy/nICgKn8aE7C48MhMFkfZ3M5dbn/Ve+/Mz39u
IS97SsBU4KvdUmvvaB+eHBOZcGndzYxBuvrBaUuRHglvU13VZIlsHOP94XrXNlzEYFl5quYPITRg
DHK4ZMUaxS6ZS8wLq+n2yusZxRxKHPvIRuJDgFh1Px2m7s7I3xWP1ePpmmXXyhYlTtOxI5xPpqXk
QV9zd4Hxw72TeFnomuqgoAiiwzfGgrFCx0YoH2272FeCK7fefywWBoVuvfCqPQcph7ArHk7QaY0K
en4eHZkWZ15lt0PPrjQh7A89m5lbWHoBhsuLRbdD+cRKydYnRFNHsmkrv9sVux0Bb6K4WQ7lbg9z
TPYuG2aFPzz0bXdJtDxSTuYDA1waUk3cPZflmCBJxF7VDVDbShqyNRSaCxe8oOXavv2WmOGRShnk
HrcWPCED0FkDcsr8ZFRwLJnwyQ8qVi5pBTlWZohT0SrsvXqMIy+bEYKrtk3H73poogXqojeCdilb
cuR9w4PAUKpW3qrZZYqP5ggQ/qYtUJROiasl2K0ppZHhFo8CRizJk+8DqJPWoiZm492wzPzE0tGU
dLLIKPh517XPbIT7yrXtQBdE3pklbknMHraXqiq6EMzvML70UrBLd1GsJBG5MuHhBVvHiXOnamBL
EdyWcVhI7HiaGUjLEc/ARBGJXMyW4HK6kjImTy9dZm8wDzBHnd9NfTAoRxdKGwtvK/JzpSOGKOMS
Q4Xqu9cFBLBCUBK8IKdl73K6du60PDdc7AGiMWHbT7VtyB396FNsnoUVAJ1ZGa/PjN9hRgYc4v/8
zX7pirJ/wse/UqYwIdKP7GQi8WkoKSw/Je1qP4rWCDKQPZAXp0RiNL9ssieaE5s/dGE6jBQSbP+2
P7Ukh+gyNydy2iCXgW+aVc00Kpi2ZQW6vIigyoQSj0ZTgsxyW757GjjjInTP1+RY3klL0bxz/7KN
/nnRFoBxNZpRly0hIb6t5GaydcsJ3Cqq61zt9NV73ZMTeVePPQE/m4veut8K0rXT8sV910qjVJ40
OTMVCNbVTpLoqCYL6n8Fh0BMPmzpM+ZvQFEc7/QEEhBioLauzJxWckLFLqnw+iX2CVjZArlCCrVR
5PN2/Aij8J885wvAeKxbaXCR35Jx0XqoP7/3c3yqGgtTZYRwjvrSlvCuR81BL30jESvt2th3hKZH
YY3kdT9hMfirmRq5phCTBAIsYONPrW/c7cXZD2UW5UcwLSL8uROUh8UvhhodNHb0iLbDIRfUjPj0
qSvSrwljvAS2Io8D79Xdfg2mvOd3R6b+h9DXgl0kJrz5xd0sX++o5225bB62WnSI0ZL0wVk/MIhK
rhjwwY/9D+rdS8SS2O5Xls//PCtEDH/2SdnMUx1FkrPPpiApZe/hbqadiPKSkBAzMueiv8m+rl2l
U1lkqqGghRyycQv7XJbN0lSW+0CmdLqweRuz0XaiEu1gL4U1O6lnPUivHSHgGmAq8yfKCPVjAFW6
IyeHsthKs4pJfkhd4Dm5EhcMLV3S8wjFZPwz9kGOFdgOgzwp6SABXbpLxPRZ8hP1f5QQ/MSDYOmb
q9ymItSVrBfPUhPEvfwI4B0YbkaFzSMchDP5keRSdWQ83Y4RYW7ixcHknXvUh0u0y1L87URcqnms
P5FAP2W8NOkA/FeVFMnbx/ETb0gCnZQuS8684YNyqzecMhREtz61ZFQFg7mt1IQE2wMp1bOUez4r
Gnyh3uRebA0r6udre/u8MN7VCLy6rlz+ySRFovdDmiaTVC2IkN1BYLOrx8BurbGBR65p/5QZCc95
81Wvsw5fPLx3dIicViyXt6ZmHqZfin3iUFObF8a1t0s8NdeGZD58QF0NN5q8HW9P9t9zH6eCZjei
3wJ8h1diHA3wcYHkD3sZnC5q9onC06XHRZCxYlwBD3vJocZ+KbK9nZxtLe19K3ycQBqLaUwmN8f7
OUXhCRaopkc4vEGnzvKO2P2rVBYBoL6XGljHX2vmDiM+dE2CaU0O1M/GU9IXR+epXygf1n786XSU
7eLmZYa22Mjz+sqnsq1fN/zCH9rk1vAJwn8WlvltMOiOD9RCJNWUmCmDa8lIBcFf7Cm7v2n+wfTr
9h0jTMWbLUquLhdVm3kNQq/arATaPBmJOv+wsjo6mAtpDGA31jAhKDMWe+Chg96MYy5KN4eQtFGH
5H907991bXcEJHde5jYkFvplLp39nPkZMBE79utpAcULr/0z+FyrVxHEBeF2DsmvvAjnw6heGV9v
2K/j6lD61Wp/t+GhGmRfOt3jbn7mYwzUH6Mt2ea7mk56BOb6oMxeh3ytJbMd0tDgnCg/V1jET+nV
QGHSJH+auWxqS4MGwBSO8ImTCDzPVhBD9bGGnNQovLgtmrbS6mKcBrzBPwTpUwnW1mCuvNhQrkfH
GFrhkCEnEXUEAds52LjIYCgHjHDmWglg96W3NEdDgN9OpfzuA1Nb7fl4z2/EbB9hBBJtPjTC8KJG
XjvJZGALtuSBNQo0NFbm9Q1lJM75Yq6QsgfF0WAlbHMIN8xVfeyJtrbkFrGyBgeCg9hgC8CFwnL3
8FJHhXDIdqvu33tHihGDuiS9h/srS00gOjRkJRtF9oCNrPjgRmxJAO5EqdaZt7KyVqIQMd88hI7e
EqN1dRiRFVkGJFwqrbBx5MuWz09ZAQIbPr/EHkJAtCIJKwuujj7AMiq2N8KZPvA5KAQviEjlaB1R
koaVuNcWwl+sknEWk/AK6vO4NulQbnuf2J4JgkwokpZoSBGxMC7rWJzmQ80Tc02ylRL5QCdvXYBr
OSK7+QCagZ+WJpGOYdvgILzvgd95/LQEbxw/IhnUl952wDGXdIfJViiynrgy8piiZKk6nWkm3h0x
ngJop6LgAxadisxFZmR6YZIOTFAGC1E1PJRdjz6zuA6hAOjiRx203AD4VxcLrqZGiPGNuep0f92q
B3nXylub5GRp05J41+d1hcuVTzn6AmJDN7bUVMCfFTtWL7iQQWRrzgehtGy1kA7eFXO2Cw1LHnr4
c4k672ZxMm88yOtHZQTvUCQASaMVRY8eQnvsjC03h/txrM7zi26XPNL6TleBMw+PMyjkVqHJHoLC
gbUS0mf3Hxa+Eer/wzPF+g1KsCUmR+vLYxZc4bEVNNGyKBpsk0vCGc7jJBRLKyqv6LO6hzgapTua
gYYS6kj6laom0n9TooK2lyZloGu4nSNx4BspvxpS6A5Vaq0hZEp9HNhmD/u/JXi0BdNsbdg1n13d
1Q67jAoFJ3L8aI6KmWp8Mj3UN1h2Un1yT3DgWP64tA+Jc9kg0UPJWbBMC+dYMycmPV8TdoKzD+DB
042lDY5dqGMhCXQgyxayRugH0GaDxWKUKuwoRLYAyh0umSFLPQ3hJYmOZurXlPZe/pQrQv6pqpPc
Nn7QuLzaTnvceQpy/aZaDCPaPFEV5AlCVwNM/RQCbT7LmWCpK5/TTD7QPCnz6CTt72cE3VT+YHU9
M+rzX5NVoXjW5Jcl2OecPuGu+nmAZZ2HjJUsVEG8s1gStJHUYK8SQEWxEHWDJ0pHJgInsiL6srG8
aarebA493qcINk/1rx+A0iQffEcUwP9bONzZfnirYx0WthcMzZcuJTStSR6n6EwjN6DiMUG6Gr/f
nviMrQI4CyGqFvgvPh7kU8VIwgqfRDpE1v8rDNZSU61cVivFocukVm/JeZ6ppebWTh58zqd0XmUG
Po3M7yKlLCP+K6rClVpx225T5fPQxohd0LrEjiBTWvryd5xMzmb975GMCU+Zhda5hlHkJ37KTm/B
lGBxcGpSOR0lq5UJktlalwa7c2PcbwHha9Ad6g52C7L0JmRZ1tuxYbMxHsc18KIOf7brx55PeP6F
Z/dDW8w2ddaWzYJUO9lxSOglp6k9u8qo/aLf7DmCjR/XwPsdgTrdt8Tgs/fWG3aHVRckIpUVSeib
uSCJsBedlw0NH5ozM1G+i8/aF2exnx32XH9XcdfGh+10KjkK+ecvukC5pTrNub7D0fz+gcZ0Rjen
5kFAViq+kvhpOdyUabyrCi1fznVgvl+S3AHl/n/iFB53/DGZpKxt3Nta5FaI3l0UF6aDA3kDqOO5
cp18tTPzQ0RrJ01fs1abuSprq5wX0xnjABvZLRStEFVP3Sb1lGJ0hY/wAK+UXZhc4OlD2DHqRPCV
okBnljCGpzJCtx9f6wnd1UInE7dKX03HCxb0An1K1cX4+TXraHfXjEYdZdd53VhVNIFhGLnSDzG0
D84NQWqSog/DTnZIB36WgPNXKlbfiHcYX2KKHn0p7hvKkoZFIevb4WsJMc1SADyOGS2S+gMCH+Xv
E/TpGeUyBdD4F64lLiTz/gDqVtMuRnykjLYSoaRhE0AKMfB5ihIsQUZfWaMG8O/BoWwculV6xFBG
S6l3D54v77HfNir/m/Yn90nOQ0nnrVGvDHainVPPr57ywJ3st6HTB7wp5izglBd4ZvgwApjdAWfv
vgpLqjK56ml5cpBgnZ4zQQ8nfhYLR96UvA24psdAH+R38lXtMJdlC1kXQ7o5/P6qL1+O96w92w7K
ntol0b8Om8J8ea2162L0cLCB5gbYrma5ZNmPKWOH8rmRxTYNqxyhRIHoLVdBiX28RPgOyRYwd/pj
MPqDWnffX3kSDJWdgvIGkkNhqbFCtfdFnrvBGbkou2Jhos/vVDEUMhAaaIgJDM03pXmcL+QX5ZsJ
DEdYNudkW5DsdTmuW0cDcptQGAzbwXEJFGMlOWSa4YiIraYR4IxwLMdcA1OR8kSLXzmTwqe5hFDE
2LJhCHVAgcNZbkZBmALbtRdQ7CGTsVNIVBhLuPWpb2s6fDdsJc3ZZbbcxjUme5SU+Lae0BLq043H
vtzV5uxkqkg+Tq7321mwrD72EIXE7JuHcLGRZ+7jC8CKm9gCLf/m8mPlDCbFYMG6KpEUJzpOr0X0
gdIAk6v0rRdLemWz4H6QsfWcO1LKNHo87gZATmY9X8T1DOMAAvHHMZRvbL97Gu9ybfiM/Hlv1EWN
EAgK2QUsCjAcSElpteK6bUM3HZalVUZqvI8lnV0KWRI/ZjzsPGRHtPpokRAtI7e3TE4tt8kvXhpO
KZI1GbXJatbotbQohlQaeHplF934G5sAeGys2c12AVHTR3V/Ll0LWBQntE/bV/cFLJCjvPkAeRTb
cWF5k14SkGjbpcZNU+uFm4srDrjK5iUxomlTBPQJ7Jsy8sK4UWRrt7DyULrfXa4ziuR9gb1I5Mxt
m9PLHSYAl2HxCTdqnpVmvQoxKXjYCLpT0hIbNFdxBHImPOckag0mHo8lORVpIeNoUwyE3bEDWj50
ESWU/KTfIj7KrbE+U7PwgAjx8dt0/tOdWBk27BoNv6S6GcZH/URU/4mEnAswQ1UhDobQVJUG9siP
VWP23THOQ7qpNIsIAc8AvpLQI13w52y3/X6ph1SlwqtxF/xU5AJMOr23ylUR3HprQLZHPUmFS6Dz
u1mX0vzcG+QW9XDwbFm/j6ax2iMDv4O83OPiK5K4s/MSiMzcK2P/e0/GBQT1SP6fw37KsCohfCJl
mI+CswosZ6GiN35/KXDEfguv5qvhurO6AgwU0xixuH0tWOu6ZF4W7ryXxPluaO0saxdSfLaUDW5z
ihqECRo0zGu3imUjyglWaqWuzujgvqJJLS+Ch/RvZqxvWgQ+SX/4MNMsd5WlW8leOPAq8a7cZFfK
gmn4iWnQT0/ak0aEExR0rAoqTWUl0jttEpAKLp3OCY29m9VUJ9tIyAgnmiQjM5m4fpVm4foAWe63
jXRBpyP90IvnwTc39iO1enuxSygg0aT0Gq2vjt5NFnJSKO+wLMRTGcBqJOQh3msgkotgryNKBz17
6XRAcBnVwGrXeVQ436CPqQpTr91A9tAWSkqhd0mmQbF9qlnlAzBLTH10LkOO25ZvRPyuCSK0phN7
R0MWqeqYC3GuFakZg4DEHmDBm0Rq1VOFNWlD7Sq7aE/3I1NLbk0rYgnYRG6To56+oPeLJ82FMj/O
9I7ZmvE6OxJsrO6E37fxaIp34BHR7+znwHmbxMJHcJji6bE+6vFDQBvgnVCcZoJWF0d6bVC4Exnv
aHrMiEe4Uvgzgz7NS/8pNfa41RZZ6GHH3HR6kU0Jl+JRCl/jzfdWjKyLmD3sH79cCJjbN4UO825o
Rb9VhvCuh6mlvjeHrQ3eqFj5Qvx9nfzCke4m6eE6fE0koMHjnZ8HIgU5n1CCyCLVDyBHdHmPOq15
JHfTUnqp+UPEQNO17dM3yxAEJlLiKqo9oari/G0syQL9Gf2iofRt3CtAqzk0CAYBXml/HdX244YP
ts7ad2zqbtGw2Rv6NglvozIhzDWp5tUcz0amZGvLnbk0JXWX8euRJo8rg+5A56n8/QZIcLGg+UtQ
PtWaiWlPHwafDzEi/2l9S8W5KRBo7KRoTkZSu3LwaeOawuMRiX24pE1THtnFioXaJC8HZyd/vd+T
o7y47Kd+4/rJf9D5hOBfvt4MCdtB/jseBcMlEMdg4wMflGLg5L6cZ0QLaPt4AYqvHxYBGpHN7COB
00kSc1N6UibAEgTVS9PtP+D8L3zkgPUH2M1z3/IE+U0jNDQR/9VMJ2oexJdgbbRJHiepBCKoArRO
y1LwyhjPOFPAeWXiILci1wYnXAYVBhxXpv5ONHZcs/ajMKzAzagWAeOrbyXD2p20LDHbvWp0prDt
JcXkbhnAnjcyvlrOJ6XgmVTN75IAjpoSp9t1erPEOeY1uIPB3ACGJ4U07+VMyP3cUSMl5NCcQsDn
ZwZIl12nnqoRcESX7DwlQmuLQCRFFAkPjt33MGGIPH5Uru8gRTqrXJGsn4Plr2b6Oovcf4ir8Hbi
GdrbOA1mJaA7XxA6iniUZjfyQ3ad+HEaoSnO1RDZXY/fih5V8kdpMyDiID7q+LFlv6y7Jg6CplGi
FWVuBDFQdcjW1w4XiglVA83p6ahIqbmnyDZ+ygUENs4McMUM2SM390vhDEC755cwZDPlnW5EqAq6
00SxMKxMecY8PiAcxVkBLmvCgAcKMNnreH0hbQG/yhlLcrp2To1BxvGomFJz1+q1LWEyg/IWH4iq
kLFEWxmJELH83KvVKnqPsga/5swMmitXOF8qbjvIoRZOG5YzU/eMtW/YV6K7bRDt8y4RrJVnQqkw
3xS0YEtCvjduYPlMjnymnHLXrp9VutBu6RJYnUMox0O+Esfb1CbCMMW172KfeyGxbJGmDV4Wmget
yJEL2EtIHJYnwxhpiFUgYn6WcmGCflbqehm4xjnm674cNymtQbFlgWdnhtRModJ74ATUfFcssEe4
/WgCAZgN8liOvwN1tzQ/5iUKDIpvWX61oIa8lXr7esdhaoeVCk8yy6JNBoV5hN1htz97F+6kKxsq
SOSwQsG1qJdr0ya8dD68Spy3gTSiULnuLMbrOX7O8sAaYo9Yfax+7LmyNFh6U0Xzy9gubF7fN1Hk
SiSh0jtnRPn2eloldctOxHhGS9iTwYvEF/nRm+ahjzA2orR8HtT0EaNv6/xnqiQqdsdBHI7xGhaU
zm4kHcDjQPB9Fdn3qeRI4Arz2f/3cnF+infvNf9Do9EZU3phO7EmUoNlpFI5tkjA9PVc08ZqOsIk
4NZkAWUoIJ0g840r+4xXv+EGSwxWfchkRpwI3DScH2j8bNVDhK8gzquS9dhU4Ln3va969Vw/6j5U
lrWdkPW2aHFbdhHb3PxelvTL9UEZhgUxt+3R40/fJZKx0b4u2CrvTZcWdNRhiRxddCOqcqKdBb3U
Jq+Q+ICI+LjEezP9Zlbimac7Lc3cm5fH0dL+ifwWtRK5M6CQm4UVTLUs4SHCtnnp6ccBM/cZBJ+B
xrRxkgPMk/M+qpMwoqCGzR3MFSPvHuigyzeDN0ZairYUdodxvPQ52kY6kpGTTbZ3p9sMeNAbFWOd
36slRuQ/JWUoypqotFcFW7Cv79NwfAYKJkbUGLRh0NsXdRjB07q5g8ly/gnDevs/hcJ7JYyhjFaz
ZrRmGrz1Hop8dF/nu4RDRVLZd7B2o1EYdqVD8l7JjgvdwYG5NKJEgvIgMkqDZclL5jgkygqzrvWc
hc8LBofXS3E3sG/Fk+o21xaMItM3AXaI6mtk0yIYTnkarWG/trOIZe97MC3FUXPZYqTB1dadqNHV
4oRt/YEBgjsLJJx/ORNt2GJJDMFKHnoZ1J3qn4vi7Fc65xZpJJ9ZTNXg4QhMtPtomk1GMN5b2teu
38199Ym8vXbJw8rnO3KXE3B1qaindHVVddDWSkWzB8h4eUlHXB4jPY/oit9DF0efUKJ6Kv0571PD
6l0GmsEbUXQa1d+aDlfexauAHyM8NhTfeYXrhVugP4124/pBXuSNTMs2ayjV+uiTaOL1qjN1MbA2
xAo1ApAziXOOy9LTdeeF3a68FN04IF6EgZ0QV0PLcyCwY5s23If2yMqH3Bgdu2+DemyDMnIaSJWw
a2S5pMWh76Ww5edO0VG2iDpDj3jnifWR/1Mepshq++XVTBN1K4yIGHNsFvYA6icBAHCDXINiLfzi
QPnuzMKGoO4fs25KONncUDTGE00V8F8Usx0s3FIpZmtcL++OEN4p6rCApYYoObAPYUKl1abGk69L
F5PoCqD//HtsaXR+jtyBh2n6fW1j80l1MDX8LeUstGtcMShcy3QZoLttieVi9ow/HDD/e6zi1iz+
IAxAnqqfmlFPlqh8nCiknpToH7iXIIqACsPMym0nWieWCrvHtd+BqbEZSpmgH9jHtYPv/b2i355C
6jHei1s5yB/Ymt7sd/VUTkyh0yZBX1/pfXmLUFK+9x4fdImvmDMmm2xRpLR3PtajGPHKurEQvc5A
TgOeRTtxzWj9lKMi2RxlYyli0yagB1dhHjtZ4qb8eQpMxQAFB3s8M8ieWnYCXZCqp2lczkiUC1eO
hunOMsS1aOw1dtF9we11wIGjUM1MOkGtwZ4Esviff/ZR5WqSJIEvF4lOktQxqf/YSBfmBOcL5T28
BGJ7vW9VOqRDALpjPJcbaRc41g8WYTrq3LkYTT4cbWNxYT9yd08pTKVed7hMwRB+C099CJsKGRi6
/z6TvSEWbmVB8RATtfwxObSfjb46A9WvAHcvC0zzbN+BhsrNDFTi9Fn87DTpDxqT4asABX0e8h3W
80z/NYZecijy1203hThVxIVaGbeRATPIVLQ17fTjtasc+rlo4FYOQn255LedObt8xdDqP6a1J6sP
r+XdHgOmRnduuwtHepnXblBzDFUQzWbQXaN9qF6ol448DsK8qOYnIEaVsWDIwzsOGnEZj8Xcy6ET
gpzm1Yi5n2uJFlf7WPxABwPcplOmfH7Td7eopHe6wHM+uG6zgdQXJaWqREZCJAEkSIWH1GJ/NaCt
PiIUDn/7E5SHPPSWJ1+zU1W+pc1Vm3WCbXAwJ0JYmGxnXrGEOEhtNUpW3aEerwa+bFvZJwDluZ6K
NlpgM2qFeYnD5m0iVnCEt2ZBs7BkNcoy5x/GY2oQt4KcYog9cuHu3zwDrhk9FsOs0hc38+5T3pW5
8DFxwea94idmuNonZa3WOZaRbwRpMtPbYPBB8nGqkLKT7mwnQ03EsiSbvYojcQWQrJABcgzlkrum
0UTvMzq2ndrnRDdVGKLw+HZfUTfNytz1RUAohJObs5+tLcd8K5TCr4t/5G2XOZgZ8QN3NdF6SwFf
XItm6hfvTNUq9i2T+GNqS9eqeFNmyRCbHlS/hQ8By5GMjMjcYLixhtU9a49ZIM4oHrpivFr3Zh4Y
v2V5A4aSbrgUNomXTyOMWUUwobuwtdf3uq9yZPwZaxqsB0o7w6sSEyL3LFyAV6h9UACU+o9tTVom
ObEkEr3/VdHXhQ7YXb++NAwPra64H0tIIGhbk/iEpDcerk4JDiRTlUkT1ubMP16qpcGKxRTOcZI7
vhr6pg5Kg2+NrA71nyu0gSOKZ1fUXE+l+LrUZ1uRH9qqaYGAVTvLgWkSvv6lmadCqLK3HM7FHMCr
cP6arHMpMm/SGQB0TcWQ/OrzJUoOAkYAaETWQbMXeTBd0qpNXWZuED778sRqhPUG8jBcpSN7ONm+
X9zSyD7OWj3Wthjxrw1XQ+t5J5vr8ktCgbensLWSHUeQC589oq7u3wM6ZkDRDzDoEJF6XqJSWQJP
0cCdDR4R1kW7j5YcGwIBxdJ6I6I7CmeWXDDhdVwUUSYygYYWiccnKKBx4IaQ8h/tBVLH1/daFRuq
z3LrjWxSHaCLCfngapS2G5I6/kwkagNbFOjl09towXziUGSEASURIMA0E6qjrhu1nxVv/dw80yCd
zTJlwbvBcG8tpOMXBn94wHrsyTuNEymcsBhDJ6QsQclQNMeW/Fx63G4F3A5w/8NszCzCB6o3Rbgz
PuYkUOV5pai7gvIZXwXHmTeXSp6y0x+zuxXIaBLR3cUe/rLcqi2lo/Aopvz/K9kADLweBTW+f7vV
OHgKag+XlIxr0QWCT0CO5ZE/y68qbCpOilq+463TvY3hJhHNZQcE7nAJATAhVWA3Orwg+kSn2hP+
pj553anoV489b1kxNGnDkyaVlZ5BM0MlWU+WO4YhR3SYlIbaeBfVQKwDr2J/x7dbURfTG7gSp7kM
/PSwpwIO2TSvE3HPD6RwuABP3CFrSllFptLsmOLHEh8ugtKQvKYzpOqwkGeUGA5xZ6MM/BVnyrOU
ClXcz+lkn/fv8Pm4tF82iZIJlwf9ojhQ+Rw1u6slK3rX2liEFAWPrhVl58mZdV5Q4iYv1G8HLQhw
NeXmM+3IPWwoZwce3nbk6i+hFqGZJ2z7ywN/4lwQK+oBOSJ/csqMENzSY5dklzYdQ+AbQriFRwYf
Jd8AO7Ega6EHQNHJmD6xXp2iF1mbNRaPSG1KIGg6suBsqVt2n8ue4B73N/MYQiSn6r+U8eCxufgX
cs+qQ+zePpjOdnUXD4pVrPYyWj9wVFhVQBj9pJJPZyNo5gPMe9OdsYGbpr4GsI99bPDHb1IHJwg/
nWlsET0VrlQFxJ0BnHxc6klHGg6sTh/6uwCV9FeBFj9/+3hAC/enbQfdTsFBvHoY2i8WsBP6ogx/
EMzx571z3zO7mHc8Lp84b3nfH0FA9HicDSdRFElSUGh1qidzlbIB1M3Ry3muiBq8gtfL3xQI8mXb
K9l3Dd/+7jmKkrb+FuzOk1kMWS3CDU7WGymNFpmt6sCTl9NFgsg9aa/vzyNGLaYsaZlnCU4QYI0h
x81MNNUnj4b7Jsxdy1v5/Dyg0MF17bnX5m1YzfIhNmX21IvoyBIWlpxJ5pVGoCxd606bCYdO/j9Y
vYPzLphBNkttXhcEOFvVPg+2e3v2Jt5FW8G1g6tVxnmTWHatr+EuP7YetSkbSFLhEXhFyG7ZYKOr
i6zTtkMghKrq6GTEJeW5DdYgFcnyEx6VRklayT4LgUWdEbY7jGcYbufijLeohF2TepNKski2rRDN
kzsFWg3oUk+OxH8je3j/smLdeVgJleZXOyOQwSBbg61tlfp6RdamE5XP+okwBcj/LJHCwCPxx92b
oSxgYE0nMWYI6h+7acRJQqQUUmLnqfpGPDcJZOq+RM1Gi5uVc9K7+dn8UkgL/y/4X+zZ3XSsvgi5
fK6B9BnTwcvuRUPdkowkMfL6uTA9zywumJpcAx6XuPGqaGJqFXtJEkWu+PvLyNKGBk/S+a7j/bc6
SKZnORZryaNzGu5cSt4R3wrFGp1Lq632awZQCmspk/qCmt6OjsNaFJQVXwEYdJeWVTeWheANdrd/
I3hkAvGHdAZ7wiOZhp52FW5EiQrSPBHTN2W2DCHjNkB8XN1SRYbWvz4AdZAK5PHGT3+kwbM3689v
9GV5ax5J1zWtBOAlW/RBi71YrlavBvjWCSHdbn+xTiu1VbNYxOSHMabv/sA8i6NhP6KpWQZ6VHm4
UlpYC+h7rLq/asa75yiWHhkAb/SYtTSjf2McvPZbmf94vrjmCllXUhUwYNCFIUYIf8ceicb0QdB/
I4c4HZf74H8z/bV5xEOw6zDeEfiZ42WZVZaNrO9DBYc5/zm5GdD7oFN1Xut7tzblGZKMv59tNNs7
lZj7KIRSmmUSgfRcP7bSYZ14C/11O3O0Sq9xt9JODARhqR/U9f4Z4Fx4CWIZSGRjpt/JeGMMl3HD
2R1eiUby9wRCnlfjBH2Ci0cqGwFMBT1GbBkW3Vco1Wk36boj9So/LRDgo2ug3AmZSh3gXdJ3Vfrg
cUe4J8OEvfMpPuGJouuhYUwqpnWg5s1rslUDRGW5Q1hEUk249Vj/VIvS2/rGyGp10Y66+5aV32/4
ziRcQVV0aLnYKLp0iMTaVUAd71PKhOTtOvk3ZUueGxi59ZFC18UrIvkfFg5lEp7wRnYuPPROaVJY
v0qka9pmyNETVqj21kBdj7KM4lHCtBBl/rlZrhhgO7chBgyI2H/RT+kzZfOZVyqBz9TFGV+IaxNT
NmVdmpyPV3ElSR8jTgK1SJ7uOrdVbOiuui6xJU4MK8Uif60pg4pPxzbfKboq6twEYvMr3IZQUDiO
P0z78cah5TpCREJwxAHnKS8X/p1ocq6Mh1a6pYkqQFeS2uTm9WSxg8DvHfvo5ZKJzpjCQT7t8yeL
eN0lAy6IkcvWenM/nXuxYw0h+XAowAXdR5ZWv2lsVU9F8BXyAuhysv4w/ye2MgwndH95FKWwAtrv
y8AaRWuDUZtnClhbazfw79ylujCGDf4lBSR5eo8GKNpnlXvxsPI/xdqDRmM1EI9AI7b48H+sLeNY
4obXvlAlY56W+1ywXhE3Ndm7bhGBBeQiOlZnQGRDXK9grgtsZwhGHFqASITP28ksN+toN7nroSnm
MDleL+g186BWThZahcOWyNiHvgWZwo6i6gEyh4XSxM3ib6Z/iu3cOk1TA2ik7z23HkV3uMa+atb7
7QoHQOj44wEd2/QH5totRnpeTO7RE9++puQIlfzYVnb5LvjLhtAbl2UXb36/dNkzn8wMItgSGrtP
uNajswdAqAcD5poqj4Ga7Hoe2tiOV+arCLW466lLHeHzfUoH/eadoLiVyJDXY4A48Expp21pM4LA
xf72EFpD/JFFfKZ/RFEyLTzQIz2gAlEV75/UYVmRtAUNtOmdeOgBiWnm/xp2Nww9AUOzPYBkTLtv
XkwGh4d0srQvjOWHBqPfQsacRkSekQy0Ag8ujiJXGNtETaXzxpMmzcDC0YFDQVZ9DzDFWaJIsE1z
NljXh5BQn3S+AdGvTvb7LVkoHdnrX2HmUTFj1Vm62Puod9nQQKS+7iSBmVDaVpF8RSgSKlZz62Ss
spMN6rOFoOAlQWovAK4HTq3KTqo83BwDRqHC1ACFSwdxZ4YgkjrDQEZPu/vxtzf/c3nQIejCgf6t
+I/r7Qsoo+o+WSjxnmCjG4Y7yxX6q624QehRIcuTbfvv8+dvIwZEeCaYkfoMAp62NpsTtPhJ7nP4
UJGVLeXU0xfYxdIBOW/PxpSlnMJ8H/hz86WAmN0YKCf+/VYTPo2EsuU+LNZO1JbkOjA8fOXDiA1L
Igq6bSG7VEg1a0FgGnnRDaSygskpkEtt+z4S7z2356EGKJbI448/xUq5JtBKK5GSuITTu16xPvqa
8CH+nZ6S7RTn4xGapxtk19Yrbii1tUiaEn7Y8akBzkJVZ2ihfeNrc7XenUAO5XAneHlyPD1/xtdD
54y/sN4v1OgohXoaUeSttbP8utZAFm4hFoR/iezwuxsZmlJqgC7z+/KFuJv51NtjX39vl62a9US/
0FfOTlav1Vi2idGlEJb5+gHIVUBJzsUcs5vA6TfoPDqdrhznmw6SG1lTfgF55lQS8+Zy4ySYANRi
vful624jcu0/pxrpm+ZNNAucN9L+HXLnhFI9mJVjhMwtudMDbZpMHKLqeEmyc60xQJgqtV0IeAvW
Dr0JJFaprt3/frkghtVtp/6oNEZY0U7noszh2yw3vCYvqeefjh/EOfzBrZRs4q9pEFQRLtZLVASU
XAiZou7XdfA1nVQaIrAFNyvn27C29IOMoNh1J6d5pzu1q3QrDC7DR+sBIYrTjJQ5xTUwBTz4TMRV
guyoQ1Hf2hi2ArA1yY/mpweM7VCEnJ3HBesfZ79NKMR2G2a/bnjoCY9uwCSGu3swDa5c1OwZ2yQJ
Utn335iYu2PKU2D6txSmZJOUd90WJ9ZPP1FdQ0PRpXsxBG2ygyqtEDBfqC4xIB5WaZR8IwT0mo0i
bCqlws8T6ufU/5Fww+JPNOgCvS4qH8lzhXHx3OoA/lKInXnT6siU7xSwqYlgWuyRZraa7+YU7EmN
da9u56FekkNBGrT+0L/Wo5RipC3AP0cX3XOW7JXR2lUV09iiIjRvQVNPNlEWzd9g4UjsXzba/0Hq
XAO7uPRKIGDnb10O3/x5p8d5zROC+Z13PIUVXKaSyWb0DICDlAI8dryDG1BzIbYe5iSk7gZLhpAa
REqLMqTmSRkEEuwM5e3aRXnUS+8MS8QmLfj5iWiVZyEbRz8tkUjXho4m910uTcGQDd5eP0nWuLE+
MJEZJbZaUN0VzN61h+R9JCWftDquke/Eox+dOi5Xbiy3/+F714OFn/7W25pH9UYcSBwTohYarie1
rcOuHWRAkZxzoniRb33beRSWBs9KCxxwK8jS/MOC8oWosUeUHUJUgNIzjWBGNp7i1W1Ti0PnR8i6
mfXwCHrgqSKtI+IFIDI42pG9Axr/eyObwJAbwmhk1Y7P03IJPixR1/CY7CC8fEXRlmMNahR2+lak
JAzwBL5wKohhFiNa0XATpwdfKGj/2wSNigrFYk67UaWN3LWN/33NxPTuypSdOyqJqULg6fwJp6C0
a9wx54bPLMhi/IvRTfVj/8dgE1RC4PT8JtgW3Am7sgsLVVebd+aQFjj5GMBhOj/ahFcL7+ihy2aD
sYR9atQ6Qx9Ey0ngS7qqFSA2LXAxBspEm0bVkpBA8vHdP0eS6aEMxp786dcjsis3LgEbV613Ytui
A082hviiGLiZEgwZWRZN9/qSyijZK/DGihyfcD9h3hL+X+LEejNjG6VA7jGea+q5pWJhEmbvYujq
lFRuUZOqHmxD13XlOsbEja480B0nqvAahP1CI/l4cdVucISA3MxymVEFMnba1tLMgJS9JmRSbnMZ
cA61M0YWL+xYTX4P9iOSTnSLYDPI8Dr4u2T5t5NoeYXzOg/V70B4tlySrNvNU0tI3XTrO2w7/v0+
fHiZ/0mSY2mmfJx9zC+Av7r18wYdwS969vOfvd4cK/CaXbG8vaf5j0UcQj2bnz+CSCgsczzBwENN
YRHTAYH9TzTDZ75BqHz8qF6zTpNdXmS//25ZcyuTG61DsN4T7d/RW08alLeFhAMKc27aYDzKOVht
D/zHqXDkaldsSfoNNmF/xg49qhi1rU/1tIgRKx115sm+scyiXlQf7wNiUKUU+JZXfp13AYop9SUR
NhSo+2BD66f5bK3fIGnu3UpB818VWwf4Ug0NBY2LVvAcXq0dCHKcPwp6V4sFT+MjfpMjiZM/QyLq
eKsVEiAHdpbxwO8xLIDQX+pq1ZnMNzbBDtBTw+CjG0PkVWL3UMJfv/fGHI1WxRwgVOtDsLtkQ5BM
d5bsTQUVi3azABbmAZ4cfi1fRC2kcC+3LCBLjxCZ5v8Wr5TuLBKObAdm8XSOmhdxNORNaDtd3+LC
DditYRhR7yfsUapKOeH9AhX5uB3NxW2zU5TCdaht6XR3J032kqWAXpdzrEnrHncpM0Lb3T8eyXy6
Bv9ilpxLLrS6VNNAVszjbnvsDEuto5WxBVosaMxhkDCXItGRCClpW5Zs9BSUXJiOB0UMNo+fqj+3
47SbAIz8fOybUeqoWQUTg/BLiCAJQaD2LEnoICENR6Z3o6YGEABvF5ZUe30drCSRV7RXqMVGW0rJ
o4zSwIx993SpVMmmVFgRZcZtaGbI1dhZrmAP2aIz78BuRggczjm0gFS0jr0KacCQn0Pd8m4aRpyi
HMwz/re4Zl8w630GCKvaNduVmO7icSZ+8OlfnHQJYpLPUnAcYP90ButMFcvQpddFBrFNksGCg73j
/NpMLzyOWLBsE6hZbvRgHyyPwmitz1eTri+kTPWCLzzLVhJQFYW9ZQX1w04CQdR9mly+D5MyFLug
JRYEkG7Go35s4uk1YDr2pIZf2q0kKF9QsYmZtk1T0hO2HTnQCIuJOwnVn0VwvxabQqdOsrnYE7pR
CUv+3sUjtzmZ34Hy9mku2d/iAHTmnLcBSjGxFkCA0ZdjY/LbNjsYjF7JXu6mb6vUGt67GlfA6ntS
R/E4CR1eiAyK/XaP05Af2yZjSKl9ihlVeg21eY47cKkTSfTzz9R9QiozL7xxiWdOov4rTO6OPpMJ
L7VUvJQWb3F2qN5uIBPXe4JZrV/L2laNhF/X2HNL4VnvJXGVmMML0Ig8DXXkrLFAqx+vODwyblO0
OiFx0vHdgKQeyupCDG8jRzQxZ9eO5j10CpBGGu5PXrtfNwlMNMhDQWLExuAfW1/TyEBWR20NyDHW
8n4QnW57ufSFmDXf+AxW3unp0HKrvKKtVWqXFrIbwlJ/XTOT20rI2R5bRmGF9lItlakMjl50EXMB
YDpUlH3xC/kujNnPTayQ5txgySRSp4Z2QAQ//wVaY5vRdkdkHORIU2r7Cq9yRCSizm4CWw6rajSd
tclzEVqeqPkaHVVuJEB9WcdS4uUKdc73MaSfNprEW+xH1wggVJFUQOJB8mUpjCN1hO3uPiN1aPV6
6zdX4gBfNz+JmKNaKWAjIA430hmxxaYLtuH2UiKMywyaJTb347ZFtXs3vrkv5gCguLbo7Ek6QQxX
KQhVrvzBVnjeLZsn9fmVZSP1u34C/sHLZ84lYASY5pqJLxVSWzwBCe+o4oTRTqtGI3aoqaJPCqHQ
KIoNEMvNw2dCnZ4J0hXe+YicguaoOY72qNc86VPTc/yHCgW7o2Ij+n9j86RXVtYZhNBFPUAgfeAc
wzW+Xn9FEUsKaxHLuZRleZQh5BZN/89IQwNiHyWGOi2k4OCMyM+xl2c1FrV58c7L2nkqTYSvn/an
6aXtpyBLq6/i6g5p7qk7LOqzdesY5mKP15s4R554MEwdJ6MJ7ThOsPDuxeudVlOqOnro/C3tYts1
Z26wy5V9q8JX1oKCFcjVD7VtLQnQ1j1WgsYheAogwOPuoadnHHvMCmaB9UtK9Aq6eLow/EJcxNgk
W2kW5A/L/GrB6j9LDsTaNDFVmufWdynoPgvimijeeU2ZT7xY8hER7ML/fr7W228svQ5WIUx+hTen
aTsOuYfLW2O+j2yLJZzHknUfSg2i8cVWgujB0YV/ZL+ShQBteZfHTpGeDq3W+uRU3OIN1NqjrF1k
vAuYpHfVwmMM7Jms+uKhQuH1/VjKSJHcnBTmq3JunDP9uwzlIg8A5BPWWkrDlTwxPgeyHzjVaqX5
8PKKuU7RJO6YAubKYnoe6eMxHVzFO9p5hJXkiJ0M2z8aYHzNN6YEC4hQxP2TyQ5D6UHQ687H7ZqK
OJcmvbJRyuboffuMEyBFtUK5KShLps7Dxn/ZTd0+fpSgf/JfJBQPezHcns56P6/7UxG2Z1xtr/wk
5v3X54Q5kSIQMbbHV52ny/sA2BT8RCqQFzlsW1DuAe/H4+eQkthirZ4vmtsxsvODirwyUdJatQxF
Lkd4MI+V5+5WgmDcnyI2tgwQku7AbedTWI2BVEzRAM05QKe/PWQe7sVEwR0LjIx3DALSDHQLwykK
VJadABRcSeaX4NYHHhH3dDp87tUQO+U+E2mftnwcLFhERGrzmTYeUVL1sMWurWAEjdG0+Gcwh8tW
PAttZxlw9SskDkCZCij6b2tasxNYdvonR8bYTM4NDuZ8Ibuc13NQxy99s+3tAnTKpOvVr8a6u4n8
J5EVsXvHcudirOE+F8lX2b+vM5sNO8fnm5q6av4AJ3NMkQa8LTTsdbNtipx7mVeiWXtiXJJcs3es
4Evjzx26FQCgUCVcxx4WkLGHXlqJLIoEx41YXbr0DwkXz+LoiVY0j/C1atV/V65OFCQyH8m/FvJx
+gpOlUnHfaoCDfNhRpvOeTCKx21R9eTLIaGNJCLP/UVEmRmuBRqLqKJQ1b6UvzRPtMvBIKHbonOE
IKJH4bWCgOXKJ6uvqQO8MV42AaJDmj9BRM8t9G2WrUsJhjYJAgDtFZxodBIm8MagEDq5WjXVJpmj
6KlLAuPMsCBKu1mM+12VQWZO69OSbbOQ/TY2SbviOlf3uMxRNenC0Ru17860l13kBHi4nwx/piQY
rDM5rpNE8uIanciVo9ba4IaK/JRau4I99zpUJfhHZIFVYr2vhlQM5rlUVanhdvGgeQXYsceZGXTM
8uS6A7dRv5URV22lnmYfUVssAXsvf1kvtCd7+0kyG0so83nf1eq5VQo7zq02ns7vI61BKUq5XpWa
TGVFARuOQPjAgyJRbZAENh67NFrjKiNIlmS/iUS+5fUpLwlJjylSGso8AjvXvwU4UYj74FJwx1JK
NRoX5B3jc3c8laZTV7kzwu+MDQN/n+UnegHZ2M/FQxLmuR/qVbNwZdshZEgoB+G8thAWQiPcK2/d
xCNQHjdJQOcldjSnEWgxARH5gqUYMOjqjQ6yU7sHVYOS2F8VtMXai/3Rvx1HX0TuzfrSBdZ9z2iU
rf0bq6qaVjBNkdOWLuwz931AkiBskXYYMFw5hswPC1RoKQqrbUKhMBrz2U7rK2s2+U2nDXYi2+U0
vabLwOypjSzdx9XaUaloRmmHoXWB5xMi2293I2glY3iXJY7RiL18gaOTXAsXCVyXhbCL5J+Q77xd
T5hOFZD3zXkLUdARWkthIhuipZ4Ni9vyk7i6XB2iKPKf9KJhv9RS6W57P5g9CETEobJy5zCUpQ1M
bO0cSDH5X2lrwvVeyC2VPidL+OgWDc6PrVxISd580uG1AnB3fV/cQ7AB3SBhAh8wp61B9oAdhSDO
u1rkyAcZk+oq978vWtu4kRMN8H4KfA0qETDSK0jknPH2C1cqRdAm38T+S3aQBSvQQhXxHjJccOkK
i/G9vIZTXB2WmgBp58XNNRujYvsOD5VFJGquVHqwhrLR3T1PJnLOr8cYB24mXonuHuwzTfzpgL1l
Vc8BK9f8pVLk19fOgETqQuRR10i+k5vNg27FftbcXUuek1Cbg1noN6BoGSxbZxzmj7xUmjwK4wfZ
NmuMt4lgva5++bG95q2Hg6F5YiUYz0wRAzOPm567w6b9+Hp7nO4iwECMLTDgSyO+MmygXnvDZVWP
Pnp77gVQMKTzyvw8KzI+oDun7ED+2kfo9SJNr2UUREMy647kR70SuCqVCWKo17FdP3ocDhMv2R4u
5CqGtIKTsuuev+FmzGBt0tO4wXENAgvzkUkWyLA5Lgqzrqi5CbdoI3FkIsROnN/f7xxphMxPJYFW
CSgIOV6FKsz/gr8prB4NILmQikKalkKja6UwaNdMBh/J9sryNykNrA1sfEoT707rys8XbwqtOzYQ
hbtR0r8ZzAMj7piacKziUwPvtZPuI1fqlnZIP97iOMHkzlr15OX7SXPpKn5A9DgLnwYz366ctTEk
8170FRcujVzf41oxWZc5Sp79UZZdG3rtRWVwW5RTFVBCEj5q74A0GdKz81nHD7pCyTtRCp4n0ceq
HOHeTSHUv5u/sSh6Rx7yPMYTELXgw1KLPXtRUh7jjdB8kaVbOWUa9wQ4ipw5FvzXV8yF5x7UNXhP
PH3UFjHzuZzKq0t/rjFFG1euNsLx0d7M30UzglIl7iZuHtIir4jFoHIz3vyR1bg9b3qK2apn9PlW
Nej2C/j0nl6dI7a+fqIhgqhG+2GkieKQaLKolrM4hzXlgjtzS7pXUpBnaXJAR4XK9Hr+pL98OlIA
ZtjVhMpzFeLG7pgXVvgQMY/LiJYxsv0RjAVIrATJrYhEb6bg7rntcMn/pNaxu34lJkydMTrhQy9S
fl+TwN/7YQpTamLKz5f8Hmvv88U/2jjsNnFxg6DzbUNJdc+6A8dh9LLVh8ldAAXSBhAK9SYU/3EX
Cl79qzmvH26ONDugbKMqNGMqbkJHb3WSraSwd3WrbkcHyemqWk9KpM3J3zqrcd44q19Kqf5mQBaG
lMcponzZ97mI4KaJZNSZPer//Um3tEri1Pk2sSHk7EDH1ReKNV/LFcbPBCHZzsFySbDvotapTkVn
8KuCk0bi53CYXhFDfGqRY6nkwVrRTioLpHkDDd92HXW3Xt138CB3B5nfeyMoR4Jp+LsBPtIF9tyt
1EwxXUmeKlVQdECojNkdnhautReZ+b4p0s3pvoQoLElmhyA7fksD02bFbBi7PeyoZZyqDpHCRVeW
xX4x/DdWBa5XZEzb0HsxEmn5thsowHP6xBivSNp4O0H16/+/e6mRVBr6yUR1k9kN1ik3IBNysvwZ
FusSih6VLRlPFqeEnBmmC+pcNJ/LEicsONpB2abrfk7bwSyKhN8AIk3CMlkjOdNuk/mnVRtaYNA4
KGO96qtue/Zkv9gwItMRh3dKmiVz3OEph05a3VAPi2oTCsbnZc29SbnFtfKEAROVWn12RTnR19S2
skQ3nwG8dRFKpKIqk3CduYkWWzi9rwAZAUHHG9pVZHulDE8Zyc1ZhDGgCrCe6CfplhxcAB7WybFn
bSutc7KBXwLM9m587A1Wkxv8eJYWUGfYqqAuGlZPNJQsu3KJrw0yUZcIZ6bpJ78mU8TfK8z+2/Mq
pqBZCdIhVKttxk+EtMD7xnAZDcCEZGktWwZxD0x9zYOLStgPi7YfKlFmmrFbhusHN9mwZUb4TnXy
TyWrhGzL2QtXgMpAy3fZCwgFzSlhitWNoPLKaLTpf5dMy3z1xk77fLCDn/Z8+5WIV2EYpJSpM8Or
K9NqqkUXmpgNIVYZiGl0HEVYAxJxCYqZE3dKoZRp/qpafPlD4vPSuwyasqkzJWBDRv5x1gL8L5jK
hTa6wTNoj8LP9we9arnpwKkMkGlmq/b0ah0FiPGXzjkZJtKymVZoWQ43URBy98ibztqZY50nB6WW
v0OtVon0+2OrrIH9aAJRX4sefTx6a4Sa7cjlbyQWA1XLtSqPd+lXvFrmwBaIt6Q8OuPmf086IvyL
ZdTOC+Tu6rXZZm+aj69qKSfsaxGbjmYuVMORIsjvpvjmdD2ph0UqUeMYpotCCCRtWdOgV9C7uPdu
1cQ0KfIqp2TiqY2JjvGTcrp3zrOWW6zalhMkospE+3KtjXvfZRlmUERqm6W5xaGqkaZRQnZI+dnw
MkNvJtOPkYMjhBialKaRdujtMUqp+INKMZUFwIuLX1Vk5aiI8MSfwXlT2PdInT/ExLd9oMRvytQK
9qFKkSi58StNEpky035Rp3Na333xvLcoShZPHM5taTizcf3GhbPz1QsHwrhKlrJO1A0HPR5m3Gto
IWADS5gbyrCOCr8Lzh6l9QSVXm9gD/qEHHoLio7XDJCDPOJR+ONTpJNCozoYoxyUTSRd3onIBKlD
sP66r9SacNWsot9Mo7Tw6mybweWRRNF8+OURa+PgdQcT+/Rt86h3w5ZosxHzhjJ/KkEB8fyTqO3K
6HqJnLE6T+mX5c3fa0Wf9ArjuTzIBC0IoEl1ccR0Ycjv6+eAE0b7c7HuXWH9lXR6SUDblexYHufx
p6yTNFxAzf2Zudrg6wIPRAa2wJg7SpM/OJTzpayH83vDr7RuCEmTNy7ipOH5Vcx2V/ZHb1xtCFpz
oTKvK8v/DoO39vaIBIumnNg9beKA5Lq4UjHar/lCBTtNEnR1IeU0OVaJUVjOsViDE5YGjE1TDXqh
6TtJc4qYFOYbFz5piNDLu9tMnYUwYNDmnk+tujJD5zm8kac75b86wvlIh7eCyH4h/yC2o2GiaiWr
C/tOCkQVjtxI0l+JbKsohrc4Fxb4quxKSEtZ8goTCdMuPlyJZ9dbMQf/e9MDT8rtuCBBmwwAgtTp
9W6r66Gh2EJzr6y9qdpK4ezhN1PnJp0l3yAl1+10mntNEws155Ijzh2QL5ejsNeu8w++G0d3CZx9
fIrkXo+TQtbeXQl9Eda0K9AMOi89hq8KKsQyT9HU8r89qHdDiV4Cr1li/W/xcZ5airMQEQUYya/r
y4P7Cub3oko/r7BVQbL3NJyc+o88qwOU/X9rxDxR4BpeYYcGgfaWkUg8Jg+9aRmAEyhpq8ZKdo8U
/s5cZHviZaXNjEIpkYDOK/S3jYCTvSzcFxLFCbAsHHw595Wz4zAJA66m0BJgpuWSR8U0v7YtlN2z
GhHFDcaJdsX+jTJx8+HivUFhBbZBfeFqia4TEODSSM1nfwHh+3sCaOwGzL/Hba+4ZzMVDG1D3Jqv
35UcBOsBti0EjCGwzE7HlAd0hKjDnvzZYGmVNg70WpNNZA1dI2fTU4l0LoPiSEPVv2TaRs2Z37F2
ZbUH8G1bGADliB6d/RKQVmQ49sbCU3Ow8ZYv+aAcG4IqgHYnn+aWd/7Zf2VyaRZHwoHzoVBEnT2C
6IePE3qkY0dDOc5/sg6esWPFvJguVSwM36P2YDRQjNDi2aDOciWcI7USh6Ai5MoPb8URbN4pbWbK
w3l9XtwPOZz/FPxgmgCpr+HLqw7WKqkg8sDakbMGycFD+EfcufwmjPhYbZNIOdS9z5MFaWwKMRhg
Dl91hN0xY46UmJOzQktQxcLpgkcpwo4yIZbKR/ZIKu+5YKTcBO259jgjZzRdUJcLFg9dmhem3MPB
Lo+mE7/NrIL1rX90rR3CdVk80JbMVREb0+8mJHpZK+lJMH9wQUkRkiWlyj4jQ3k3cgRuc7gT6GNE
5HF9cnllwMesxvJVPX6iNFOi/XVrECvgNo4/U7aAa8jUh+GiflxRMIhd2oZEkZRzA74msIApNFk6
AnalgLn6ph4KxVn2XXm51eFepcHfuop3jgEOnTZqueMwLziBkpj6VvaawmCMohdG8OKVz9Rwxc7f
6/ILBBRt80oSz9rHrbeCXxXE2nw0HbVOpe4R6m+lMEXEnxAUodCmbXUxOuYUyKum5VUPZzx5KZxN
tSi4Bflm+8B6hcbEXcfWFOa7a7KuYwzGeuWWQfItkQlb1s2eXHzGCMcPSoBGUYDiT6Us5+HYf+ir
Gp1zbCchksIoYo2Mud27Jp4GfeKLp+btcFc141eFXmeBRfdVW4KVcnNKANRDXGzRdD4HYu55Rl3x
3ydfADhPCY8HcfB6IRtD88sXzazxprOToba825H6XyS0SaBk1GyBcyHAcLbHktfEX68XS5LfHJWf
M2P0oZZLQ9qaMiFx6VuSRA+xNaqEqjaKTksLF17wGSAuvcFNJqIKRBN32EguWsJlfgb6FOXOuGxw
rmcqAxRQ9MIftwfIs1wwzrjXkyIJ+UwhW2RDg6IsWeDJIHCPi7Nhnw8nt5T+i0cBjmPGym8vBvSR
VfinZ5cAdDG2KwU1DYgOBYE0+/9axMjeyqc4SrWqVXM0moJlBSLaahtSkNhFEfiWWu0Au5H1YC/i
zlgAxh4gyjNOW9m75+FtUpWrpOPyoTCiZHcj7+zwoq3VssTXipEjdOaXBy/e0OkhU7mU6NpRDVze
QqkxEEjZ20KIPy7xOVFzNMa9GBvIyPMcmiBy4eabZb5QZzFzwcTyiqHx/H/34L3l3ILl3KtYnP9b
u+28u3j2YLyMiMFq6CZVYZpQoxmWpcD4dFWGSImyza8PbVKAyKc2lkZ7l/IzRqMEZVDPbsikSoxs
yWP/7pDTzEjg9U6Q6RP1/yhcE/Q5Vd4UXLAp/4vI2cQtaSHH9HGUXPdLsMzlYrrJGWdxzMK5H7yI
MbhpbOIAOUULRFPjoWcCFM/p0WU0VbxDVMBU+I+Ss4UnbUoubOylF/OKJgC4/LT4WIuOQX+3WZ59
3gG3jTOmC94F6VnXPnSUkB/L3ufMXB+OYdYPgF7VQbb9THkKeXus/XsBBWiA+nkNb2Mb3NVpERZV
lqGOonZXdrrjOHmxKmg/durPG9FMbkWQd5NGrWGTFDR7jfUaUP+GJHjVUzP7OSGHuB6T+F4DN38F
7bnXbvmE8yISqltaWJ6LghGnzW8ucwpca88syOvWu5+Fw6p1C3uU3RD6HFcEOz38vs4ld599zqKC
Y+3xVQ483xROA4AfvrkLoMGxKpquc2R4qzLrd8CoJfeG0o0ga2bH7kmfW5b92tCXkuJ97X7LXFD7
xJPqLpI5evjI/nyW5Btdy3nAktrOIc6oVRLgYZMdL5wv0BHpVOnghcfKXprJO7ZjWEE1Z4eoF9sN
Ii9kB9c02ONHdH+y23vL5S3F0NFiiWCWaBB9a8dc/eoEW/508DjENB+sAl67pmruvCrBZFfI4DPn
6ZYI/48aofvc6rxMs5w2qTbuv9Mo0PROdxUkTUaJN2Qvob0yKvu92QR44Qf/tHGhODdYDgHXCmPA
6XKjp3lPgXEOFa0ZB/uwZJrWBUF/PtMH8RBVK1dO1DvBtal3rpgCQfEIdfRbkzDM2LLs9AAIYKXP
4WujIxWY8SX5IKhJVBYH3070pibw6PpbhTnkshlBlcS8R0kCCVPyHf1sbLyx8asYfh9DWp3M3R0D
Nri/PvuKe76x5shRT5Apn25jONN70ZgCkQmYLBgNPe6EIvQTs8olrB11M2jqENWaasQ4P6HuLMiS
6UNrTH7P3ouemppA71FKrPwRyPfN6Z9cJaPdAFYO2dvjUZKfSt7pvX1UD/wap9wuKfmz6GPn25rQ
MxPdPmvzDH6LEbYYtpuZM+a6udaS63JmKRfEUa5ShDb+eIO4S6WbZsBUVyB84VNpQ8ClGWsA+AJ2
bENoyoQyGuV4vnHFRdwYE+SW6iDHhTerSeC91PnvNiCyF56ixFtgVIXHKA39NPtKKo/QJQOCJxt5
n7OTzgbjCQqs2XkQiQFPhzOR9Abosiy7E9GzjcogshAAhmmR3kl4XeLnDE0Yz+qa8XJICPuHfCRO
l874MyT7Awf/pibQ5ubBDO7jn6plwnA0Es091jq1O/egBLuCscGFSHZlRuMtnRrKWsLEDdrod16l
SRpXJgYZ91UugURcFLsQJ8zvF36OcDfo94ncwNMupZxivoEbjvf9ocypGEXlaYNibU9ZZ9hm8x+a
gS+XD0fatp1lJ3hzG3giSx+pyZ5UblaV3VTvb+ozMskACvd97rBj61+s8Yw2UKjaLo7lN8F52vCG
8TEzpa1FLHhfemdvh8qgKORzxzaYUwQ7uybKYlVVIz7y0EJDrPIu1VKz8nCKDrVHvqWY7SX3ULKH
ApOfpwDLGfLktMz1HndRh9U5Vb6IdKv+ZpvIoanwjEKUcDa0IxBfD0fikVCNKZMoV2iwwGFVRwTA
k8tXo1aSFgBop630aWcOFNJu4cxpCQZ/VEWUGXEG7nHkkfVcMhhVmqmFEVqv7V6lxcDv7vMRaVA0
f9aM27QsBeslcUodoJj3M5t0qU1zBuoXML0iDz5peSRBo3d57CtvLRjBKbMsAqQjkF07dzXXYdRY
GPyLav4Xs19baYE8fF0NYsVPpop5C2X1d6/p1/AAGqFLOvmYXyIfrucRHpyuaZKYXKQpxu12+ix5
1VeYhSbdUnu60NoZBRa5wmuO7amzlKCwhAXJzRJmq+B92nYwx2FT4Bhr4pHl5/qVOL9+JOi7sUzC
GHPqMqMp/58NxNv1WYTy2NMDwraQt8jeDRIzob9ccUFcXM583k6NqqPZQdRrCsRvkb9yz2h23Fuw
SbG0HaqtZGFgYlMgIARBmQoPMLWFysGbxyqS3p0DtxgyV/ufWUAQaqfoO2zWIHO/7YCIYtY2Q10J
iHiJKqQFo4ZGzVDq3p/v+K35pxXQfQmLoY8jFI4Rzp6rAJZzN/H4Jj6efDFMjsQV/Y01HLfeFo/l
TsMuqZc+Nddp2PL3ikgB9+Xy7WXBtwk4wH2fbW5xjIngjYTgeIQuwu0AebFzr68uzyIcF/l+YBmb
JljW2pmIgPVnAMvQdtZ9BHyjsvVmnLfTwmM5kDzXJl0JnPodGYq5PSqatPD4B5MLv2BDCPrkTLP6
ktfMARecCAxZhwtfOcbQEzqJszBDqHcHyZnUVlhXVbTIoah73r9SsG1cIyoRMiHo2TTFodBR9pJ/
fLJg9FjfK9sPy+P7EocBTH1xneZmxjqtll0zTKwwS09iYOi2BlajGX5i5MoVCIom5aAIYqimIK3e
Ns4fv4SfqFe90CX1Pf2voiUDMcz6Nw0xnAELVrTzZwgvHQiF+k3Fswu8ICqz1W2yU6J9d85FXy9v
iauK2R0eChyq6xicSxW/KhZXZy7R1iCrAleZg0oxQIP3jRCbJQ84KNzqT7FU8TEpEckYd5l2knKD
iyVwyQs3IMzke0AQDLT88bXN0SsOB4rbiKw54VItFQE0D+L0EszTDHkrRCDVmFFeGP9xTDc6FI6M
U91T1iQfvu23Kh0Fp1qVjMY7ehCjujQA+I7X3t4JaRmgV2gLhuZP2pfLJzivKBEyLoiA5KtS0chA
yst0RXowfhKdoVspB59gpPVW1bzD7xJMdTXBBwstNmNt1uQVjEshED6JR7XzSZLJeKM7JY6ZOii+
Vfa2iULU7o5R/lviMKe4334djuLPpVKTAnOfpnV7rY67ZLWIlZcT3ojcB7FPTiCwXJ0xWBWGfWr3
5OuBk3AWAFWKHn8EbuBtIqFBkKzRvNubJrGdAOTg25G/2zvJoEV8zWO//j24dW94z/cp8aH3BEdt
/I8PDcqqg1d2xRWwEWBYLLtvvU6H2ndsEgEyT7jXpZHbRG4PUJkXqjnxNsgbG9GiLCWl6kdaLViz
rrBj/s+c/U3oP21fa1yOjrB+k0qNpxF8qNk4UJGfKkq78aWIwS0fcg1zu43gpBYnuZXAear6HffB
w8YzHudJ81cDDVoTY+dDywkuaYhXecHtXPp4UYoE2ug740widEnpVq1tshNMHF6+mBbbsHslSdDx
UfTErrjyFVVisWBjrPeZYetjhwlQsmge2Mp+eKTTMFsNOcRJ7hkrYANdQZkifpiWHwCMIGqilLAG
D2SuO1JiDHWXCs1YvrZGy/G5s8DW0Ri/osemylOXlld0CPDsNP8HaB5xLv/Kbv7lLN5Ed0iN8QWs
YRvZ9CByvaBpO06XvbiWR3fT2rQLr6X23k0E2hkEOqCdeTDvk9XAmR4e5gHJWvWj9dxJdFxKwmJN
JKgP4EDMUSWHAISN4o+/jY4eUWV4CgjtwkcvJQCEyEQ2rA1xhy7o04obFIojUlo6ifMyntGs/hdW
JIk+7IaMZ3BOyJPn908sOg23oYAznpSW1oQ11TvpWYIDJ+setgDkXHyVUVDfkn834jZgqhVk2GpD
w952EuuudTXIyNO27Z56nKoF347+TiVx4LqZTZSssM0NPfgm9duS2NvOFOymlapxWMqa8uBV7tBt
yXLyZ3iVyDGC5O+cRA9uTLlw3n6Y75ID+fBqgxEpB+FGszAAtw69JAxlLcfzIhEZLn3WKACOEYrc
Ifcy9JXs2OY9eXRd9/sno7lKz8iHATtzPRhGxV2UdBPB/0l1aNyiHvC41vq7mmkXDugc6+nkLqxT
R139QKS0tkhM17wzhgPClZ9IsER8TOM5ouk20WK/fyIAS8a4aedqg41+NG8ClnB8I5RgKogO60GD
ireSjaqfHy+Zmk6N+xeRDLwOj1uWm4A3QjKvtNdj9AXUvKLPRmmsSNYfh3igufWH0Qnoz36uKwjg
fFdeUINzLCu1R6VDLaStmVt4xeR8SWRRhuTW51HyweK8PUw2+ZnXDowZhPNB/+5qkFBekk6kdNBX
xfo+mMLN3EkXrU1tAGdG7M0GFw0BIY0wnxDO0nvusYM4I9rbQ1/U5M3TEctzMOAlM1KnYKoW/Gc6
Xp9TQwonms8QcfRH3LrNl0SO4EP0AFMmrPKu0SX2Hft1VJVmpnUqc0iTYzpQGm4JvtbAatrg8mv1
Hhs3+tjWBNklLtHmGueDihkhqvfRRFkynvNEktyUY2tM2zLbKhSHl2f7PfC2nXMZ/dqubLBAguT+
42b8BoF6u8goo5YL69UQUkeoWVc4GLuUHP4Gj22eU/lVA1zmBtYrnRpxd0M3/dENUKqz8HGvm68v
dPmYRRRFCNo9gennjD7Yvp2J3Dsvx8iLQm7FQvE9kWv6ajYA/ktvNk5Biar3X1trYg5gTDzXg9UF
M8HCx3UGkrcgAM3zverViBDLt3aAoKC3biVwfPOW0Iwqci2AzRUHINxmE02SgMFvXV8QR+FJa/Sk
odCPDRtxUMD1WsLNpQClWGRGSttrfGzV5+ciWNsjP/WB1bEiiW4NDMi8Q2CzB6xKL4Rte64878Zy
Wow4Pj4AiJd7dbo4wV15cShRTNXk5hvckW2J+6qgTcMTceVFNYBQ7yHxhXBBy+6hTN6RDyQkf3iR
Rqdp0PTQTT1RczJlgeeoRS16HtYSliijsQSyfKpJFp8km/Wl1AnwOeeY7QP0q4yI/MrOI0l1Dsqf
fxnaMPBJaDUBnLH/zQx4ykIkhH3b3aF96n/otw0MOAu0oHjR/0AeblULidccO/BzCHU99rq8Kado
ZnyAdyjSTw+GkIDHACUsRzi5r9LWhvLJ4pAZL/P02BwHkTAqIjv1CBvISvtigyiAnnmXyYOvvbXt
tqU/nX9ufGF24qOIJhwDSWfHqVzyZwnREmHtq3qXC3Z7IhM7BZGQNxfEHWJHZex25G89Qr5iWu0j
nBV+okTacZ4C43FHiey4/E0BczqppzIBT7ydcru6f3A1xae/qnEpfKUi3XFStBY0ttkvqohDpd0+
KtAPX/cK0tk5gwuMxiE3sUDh9+KHrlztSEbCV5WKuO5zrjfagZ8JWApWTQF2xlgAR+KDRnR6sYXF
+3lnl1pYG/6vCOAavMwUwtPXAf4/MKN2+8YUMPN4j5W8pIjUZIQtaRtMrEir0KoXCXDHV0LVM56Y
VX7l/hV9TYADhY61PEif4SoT2hK5ItbdCc1IF1fnZ0jO8UE9DtTLynYbOpNH/K90Ggbd3YIllKtu
uNJoRNAwOjzHgOXCsMzKQNv7FboMqtuUUR80koPX+4jrhjxQwjZUcWNcMip7Pdm1NiWnkEnNW4pv
3SUBH8EaHOoe2CzOcBABe2LdkKWqxqb3q2ofU1jleu8niCtPkE6+VgItlhq9w6nN2hcGzGf7/jHo
jiWq1WGohQe/QofG4F1LABu5UgFS6d1MtQNSMcumVrAyQjJwJtMtKyFT2pT+KD3SeRcYy67LJWW4
Cud+DZAbLlWfMOBOri2b21zA+fHz0hMkXEl6HVB1KPdVnT9fTix7V207qo8g/B9eIm8YCPD3oZpm
iwwHNFA17yNtK8fs1FTttKPmX0uTu7e1PoG1hCk+hno02Sq3+YS1H6vb5FBqUCjZf/nj6Sh8e4LP
4nN9DOhCifdL2YHfMGumk+v8ivHukjBizn8WOuXYiO3M+bzNxdY2ACsnpkz9bdz8Krki9557pTxc
b1+zFPNxjtsf03jH07A13Nbq0GirN6gaJkqkA1mjqw/YJSdurQft8HpO2F3Glx4rS2Jo9PMPkdQw
gVzMV94eVaqJtnGYw30oIueU4FiLEmshY2HJjZnk2jgIxGCLaS5h7WF2Umxt5bHA5sPvwH2qBZfp
zDHidjhszMQzTvGjQWraAEsFwfMpUuFH5DI81whvlkpeW8/URteqm4jqbdI3pyYegiP4Q9GD5Hbk
3tFYoigacUyN20XkMEzAVYThfFTyVAW0j+sdCFFfOzsrDVvMwurOnmudJFAQ+JRXttBGh3WJUit5
WgVka7IeAvpsUsSOh07QSFqrgK1S54ThCcv9V+5npFQ9/XAWIabglRoXA3BTbGr8x/3YSmamCDve
u8fG2T8oSWtjK2DFsX5mw6pB/gBEdu98eQB5xJrH67UBnEyEgMyFk0qgIMTG/JqT93EUO2k3/PFW
co1IpvpNFPIvhV/TUVbNquR1SA1lMiB9yKMRk4c89LftSDURXei3AoVUaUgM005C5ExvV3Vp6eBA
RWfgH1au48EyeK9jpsGIA5CJM7PYSZsM6v2KTB5ipTstcKaq5R52dKpam4Jmsg0w7+47Qs3VPAsO
178iNAIJZ6wm0emUCSyV1pOR2+fWXPpfMBYktr7DhZdemOnaHaac3x27F/dxH71wL5fZP9qQw0ce
KI6I16d374YhXyPDHDiQ9SDgOig6Ws2jggbSxnEXMnA3unRercawaEunP40rxybGrjXE1in2fZso
1IcMmR6Qe4Wrm6j/iu4D2SF4d1jWerWmKgkzo91pedTH9bIjrMVYLwkSIQ6b9SWTWpIH1as7tZv1
qqoT4n+IevixKbF0anP8ITJkPNy+WT+8LNfxx+raCunYbJBjFjCjjSwbqcK8fO22yoXU4HEActMM
qcKq3cy+nsv51oxrWy/M+d25R/QZ2kcRQq3umpp5Bz/btSzzkZhAqMOOT8DGEiFe14ZtvWB0XvF+
zchc5agEcTK3kYBuzkbLb01eZLucJKjkhle/i5fbBi138j0BB7g9NdKLFtWWHHkQKsfOEZs+D43F
zYSREatUHk5XVuZmx43p3fD87HcE2WSlComDsCgQyAoNlDtEkCi3ge0vAFh5DOvl3FqFgqcNuVas
CIw18lJ3efwPdgKt3XrHx1QHyCAurvYeFhvS+VfXxvWNv7i4QU2vq7KgUhxTsy6mS/AtqOi/GvRq
p94N3uZidM8Mcl1m3O6QG9e1DnGNgLyg4fYyu9HFYxK03zmajEdgh6pZgOlGzYTVcMZ+p4UBQeDg
U76Fk7eGKn1Rq0B1/zHKrcRciI/MXnzBLXsxSkMly3IO42iWr2sKRXcYXxUdudRRm5kfPNRQfrt4
aicC5/f1zEA2OUuIoqHiO66NespzWAdNsNANweQWfXN4ARKbGL5mogdgREXxLWs3oBYDfL5CKzE2
xr+ba4Qkj1HyLNikuMszAg7iFnQLcy3KQ3XPIBb8fl5yXZBL5oHmSWpUUfe91A82SD3V1QStNVeN
xTHiF8Nwb6UT6Py+PeixTdtiyjuVwllQX2o4bx5NRd1Wxzs6wMvDd0hQFQvZ5jnugnyfGG8K17K1
rk72YmLDGE5OU9tGHAbcXSBRRwhXCtVWo2DRlon9IKrnbbfOnyYHawNOm2Dy+YLZf0Tv8KVt9qz0
9OfABVOfUO6fPdOnCawKCzLEJwzkDe57zDG2RTNd+87m90ghx+XGdh+D8utOyQEZgc4H9jYojXje
RzBEtnzHrK3k3jV3N6wYj6pNCJjKrW9nXqv5TGKt1l2zI0coJtC7HWx/Ml2X3HbbcNwiJFNflmiE
Hl/TsrdHfRSiKeeiACm4gepTdFEAlY4uG4/qGU2B4kSmVQ2ZSB4r4+cvCPt1ppIX8Vn6uhpjEfm9
4QusFneTRmZK6rR34D0IrZTRT1cj2+iwgFFJLzKifjqIAPJYxffWAjNFqtl/lmw6q4SFFmw8BJWO
KUpsHSkp7rjDLbJz+uBGfdZ0cG6DzCB/2aI5H0BbMFuvzgCMWL/+r/5xjcSUIFImvWjFr1v42Ghk
nkQQJouNMMGE1Hkwp4cDqMijLzkDmKAxJ0L3DMVNL8QTvuqzm/HwhoJ604/V/r+rZCBxIRIxtwxg
02EBQkzaB/ffdMHxZ8kiIIsg0nfBoQAW2Q2u9DjTafXHQPoIS9IM71kY64f86qMRj4gRd/EYnaYw
oNqlowtHFUBHQe4l0M7DrclBjhNf5lFXKZhGwJFCBBvh6RbHMalMJx37PTLozNBmBsAzuH4jfpdY
DnbFEusuTrchToUK9hNZcNc16VyjGhepxdiz71Lp8a7PIwn6Kve61zrvE8whc0f+iv7yobAGcw+H
bm96W9vLP9ubRcSbfAFMKzqgPj/PTiXONyk6AqcLmVE8RsK49qFiHkIPTH1yca71CHMrscSwD6Ys
uz4HpMsRLyp1fZbEe234L4NMGY7+x7kldr2K5iNCeSo4UsWde+RsaNzs72ZN+EZZ59xCLiLC5uc/
JlmLU+MR6Kstj2n7YsuWfF9ekFEHIFztOeX84/zgfcqPymCh77VI1AOQfRppgUDuPpylZx1s/M1u
a+a7SGosBzC9Tt9G9X/ufSzRbDytNnmUU5e8DJ3Z3893X6gbFGYkdOdatuqRy62n7lFIsBG9cc6l
WcYG4ABnlPQsAqmSoHznylztkwblJ4CG5nSRJYrmuZ/Y7M3X2lwWGQOs8nVHwdRSvlIHX03DhcXm
mOnddHFxfa50Fut1gcRrbogA/BduNYRrZK/e14FLL8OB30vOuWRSW9A0Vt7yV+hhQsJ6tF86PA9e
tpj4hDPeEJUrMAIjjcIaNCErsh9COJ7JEKjKn4OsL54KzaYSObsn+5gNnNIvQODChjIF9UKT9/5q
zynFvFUIptHEL5mKT6/UEusAhXIDa2Iug3sdjLA8/26nrUwuEipFznZATs/kjmoAyi6SeRNT1vrB
/pW4VnbtD0t4CecKDSjOU9tAmHwgmWUR5P2qWBrAfZZ5V5ManPaeUVvSfC9tb8GRvC7Tc2SnR4Cg
0Ho3Gazhww1EwAflTVKLlRFh0yeOjf3oNoDyHnrcTohSe1GIxUPWSRxRm7hIAyC2AojpPzMogde6
C4E3vdKTAJVhm+N3ItQoujzFGszjjQybze7EEbnRkwzjx2zcStXf1Mb6Ab2mANTyJGU++3YoSVq/
WhuDIqCMHhP5yYdGGRctFSS9EIjcPZB4gASgOlKA+fpznYGzuQR0dQe+rBWHdgdV+bbQb6ne8+5V
BR8UsQL0kzMBEt/c7cUfBx/QWnPK3GeJFSuGO/DVbHS8xy5xtwqG5wBauXdi6s+C4IcBDtnKPu4+
5y6bPSZDw+ss2MxqGCNXPB2qUGVFoyxg5H1qWpm8BFpbSBD1+kVwaz5Q8BEDWfIJ6AjmERem6Jg6
5t8h9XJUEYJMJa/BanXw0IJOVtWPz3+ZYN1SbRWqszbpZmgKx9LZR/fcvFPI6f3vioIGfrfdFwdd
EYa22bip5oKbOTv8gcmi79rWS1QavQP4VVzbbyQvX8PMDU0yId1adauOz8KGMQWL4zFQg4BKP7Sw
gjxchE6xrz8wugfnkYulYmjoxreVQcP1qir0Ii/BxQo99qA9yEtF3JnlOUOgfljN2ccsrC6NsViJ
nC+yP88iKY68gzb+15ZqxhIESLJIbQvtNirIge6VilDMJZM6/lxpXDraVREewsdL7ymawsyUS8jf
Q2Uk/ozqBAAMt7wg6JXNPiqlZO9/QP5zWCJiAS7lv1Fi20a5mxsvhxt/DNJTQJnb7OgdS53ceMXl
5380gMEDQ92SxV0gGITiC/FiSrfsQJisWUJy33rzXW0+cEUC4M9c1w+7I1dPYsqbmhXjVX/M2nc8
mBdeaul8CCpVJ1V52dRswu/ggPT+Uo7/Nj2NEDvwsU5s5NSqLqoG14OnbqiG5RIDd5+15I4LruET
Nk+SdQlpa8ROzrZqjUO7TTWwIsEy66w4pZFC4tbrnTQsgKi5JVnLuxQD0Hyp9mhd3az5/Xvb/sGj
ca7TRIgnaWOu30w9YqS07gSGbSVpRafhdJqKRPeBB3l87kahijbTKn2rqWKYEfIgLCyFV9h7AmFQ
hjkJCWEXeuZca6ruSy4tUJ8UOCuwweuawrHo3pMaYPODVDAeAh3zNiRCtyPpWvHZt/1KK8rEjGi4
lmj/ZyhGcvUiD6/1No/QzZxT4DA7GDg/RBFGlP8BlRVt+wH8kujN/2XV3XcAfxkgfx3vFWxIIy8W
tTWCV36qniw8tduTIQVLEomtQ/mnwm0XXavKLGTYxBNnEQ8wverfvhIy2n2+ntoyqiFVCRSAwMj+
rQNzKUa8OLdzh+saLHXfUTC5qy4VmNyH7SAWvbVy2DBjKKUABYXeNrggcr5iBcgV4GspShnse4My
z56iO0B8N5d0SSndibtrbEHKHokFigdG/ukhHbMPzoDlnMX8x4Av/dVcLWUv4jVogF+4r4wO4//o
MV9dowgQ6pTseCiHGDOpz/AAIXbPif+L8B4GpJOH/i2K8vfPnAXi+I6fifdLMMXFFFApsBoR2tz/
acpJmmDpTPTvGgdT4X90moEqaQPPjw8RqNKhmH6CB+4Zk17DN7ioLRpzkgHiPzzqjT/WPekDk1qm
UL/JRJCmc7uhtsRdilg/+YkneMtLlzLN06T8Q2DuLloEqO6pJk3/XOzPfMo3HN1XeNowrU8LxkJG
lE66cR7Styt5lB5F0OLZJv/aXVaMMvnWxSrGwIMPvWR1W1aEpCL37sm4LKNe+b85SLAwMbVYojEX
uno3NdpWrSW9wd1VzO4fDaFWQJ2SddkxaDRkNWYU0HjrFpFMumpYXAvM8/iFjh+gdUlAHMjwatj9
Wwp3U8fzOcr1J6itnWHUC4ZgKiPaR5De2vTZ5Aoy91mZHLOjzXMINI5KMVb7GBygXqg0+ArbkuW6
yzFLevj1A28JkbZiW8GUTJ0PMnAHdNerAoA0oADWsNtO3QU8PZooFIOrmaE3/Uh5B5mxye+qx+z8
BWO6p9dGg270uv4bbvtp2CTC+AJYxxZr198uD48HtQrYqx+1sslXFUJFB3i0udwSRZmXAfEriNxm
KkJT4naivNljlk8qC70IThNIPGfyV/lzLsSL4ao1no++d7CGiVztSjjjjvW2TkWHer1V6LPhhui9
m7U6jVqYPCHFkr54S1QmBGB1X18gIYk9ox5oSPh7UEJwYrQBCB37+tkV/KorVcvLH0TsUZ/0encz
3WcSP3l0HRPbCbyEmuZOtBCyRXNZU2CBqae9EDutmVnFacHbeecd7g8oFKDfcBdq6Y31X6psMfNm
p63lb0G8JzKQk6Z6xgBg76oDjYmxGCaHA0snTgeZOFI3KKntkMqO+tpShiswb5pRQq1B1D8cLGbG
sdf3jgD//OiwTTk+MqnYUXo2MHVVP9cK7Gr4nHZZwjFoSxTSN4rupQQOKM80UFuHhwfbkVew08aC
cb5llIHHndAveScNXE4Q1laWqFqUBFfHCogG6RNMlESEtNus3cGfnbNqtAafo43aGG/wFxG6C3Mr
7wPkI+XmOt1N2fDaNMMHrq36RfAH6/EGA3LbVJWintGTqKDHqkF/aZulu0uBMJ2i1KiCwrkkKxKV
stBxR6Xmo/F/dx10hiXMrGtcqbVGgJLM+/VCGg6tFlCs9iBJKOiSPAIhr1cWLRb2aiErUw5odXEJ
6VXGMhqnPTwIxjnMmDimFheksx99DlVPKuSOLAuSOb+8W8JL6onPoNrE0uh5pSoLtggfqwjaguVH
5msaEdp9lJ1HoSjXxu/wITY1TSjfKYC8+1zSdYtzPmXwW8bKTI4EkOjX6n5G+9E7tMN/er1Ciscx
nf6WKzchVQeiHJwM2f3+DxW7MJK/EaHTbW1/0/S9xdWycboDOWzTGzTvZ6G7Cj5bPoBjj71qTijD
cZo7ogGAShl1ZkNItB+499PZJXhMKZ/Ew2tF6DfLprrZqP+yJ2XeRY6JfonMk/1b1yyGr649MRUD
7N67BPzOtR3Zk3Daq1s+IHkxCW0XHKv2xok9+BwKPBHEYbrxDbsH78HSmbQdYjml3jybaSr9VkfF
wkTyPIPni03DNeXhxLDbN66ki5r3SEJmE5Pa5h0676EbOI8R/N+tmQamWmSAtQKjM6BfUE6o/XPU
IvZqXe5FSJuEErH2tAoc4HWjmbxAIteTFtgUz4T8CD8GmA6sAvYcdbH0tWY/tysRIL1vtL4dAibb
WvF+oYYJQaDP7vIFhFS0JWbSWUrqiv36YIUirpnGQcOrTntbt/mpwngoHCqOdUbZ893l+SS66X5b
Tjx4qCE1KzUEoa9qkrViNu0kFl/VaOObPPsqV9SArPJDudiQMum+OyKHKnotS3PU2/QQV0NMY6BU
gshxmMm2LQ9vgvCK34pWzIJsRtColoI5zfU2QFo9Zw9rBtfZrkMDJf1uLqufkmQpEl56lmUY8hRk
Y45xH2o6iIq8bLb0ivJlD14b9EEWbGck422TqpbHXmCg5khod/AYHRe6vARButHf9r+4GRRyL6eR
b00qVSdeNT3THRxrtlHUYOIPUXJGlF8Rd5kqXGQHBOGcwSO0qFP6DXNT3zbhiaawQse6IuTmDbA+
QTL/CT0rpbx9C9wNTBFxdkAJOOXqr891DWC50J49TrNsyufA891divyyfcEo2zHcM2ZFWFtg2iQ7
WTjhtg0HLvbRM8PnT8h4PzY3bEGSWL0vzd4VWcKcRdqGm9FEkfH+qEL4kA7C+r4uFcQsa5nZ42+M
TvnVikZrOeOl5UbrM86CLQjHWQIFy8EQg9KuYDMmZX4C6OE7BeQg8+22zJf1i/MmTjRb61QcKksO
BtDjDdCevlJOkXBAMF2tnfM6a1ekgMJpx81dnYPm2jWo9rOcCSYIc9vSPRGOK4uoYZql6Jckn5kd
JxfONHoR/lSho3ypyHrhn5H79LX1/+8MccyEEimTyEfQvpZKTm0FmT4e1Cl4uwWA+SauH/C0nAJo
kCNY70T8RCZeNMlwYSp0awIRvf07fznJ38W+lxGBEV4uPhRIgdutaSUOZaz+o5SAXdgr3vQytuTQ
xNNN1v3P4V6LyPEl/vKSjCyfp66VwbxXmwatWgfToW1FFBO2q4ImixJChgPaK96T8RJnOtIgCQQa
gQ2U5R99e6XX6YEgkLLRh5UdkiOrrdzU429ehEhwhsTJzmDRIA6/ANkhAFUG7tz5lzBJKMwpveLs
Tw41XONhWmyxDsr8OIwW2g/rPlHvQuas+/oxgMunVotI2xhbgflfhZR+1tvcAH77TN9DtSiLhxmW
XrLSiX60XxatfNxfBTyheCeBYA1JSrNdwYpx24wV05DcQcQtWu90AcYheHM082V9NpqKr+z1Gp86
NK70kuP92bMNoOFaHMm2KSfE2dpyozIdZ2YkMPkzd4tIXZ8Q5L6Bw2BVCgG7iGu77aVk1z8v09uj
USOybwgzpHyozP4IlxxtNBTUAyqwT2AefKSJMagAmXlkgXF92p+Anrv8ahHsEPRqrCVNEI/y6EZ3
T3Kch9vklK55d84S6HsT1DX1RvMSzch7bKPB+xNewv/+/ACDCVpBz0kRgaGdcPJkk5z3hGl+yyyA
o8nr/+Jjzfku94EvHmtLIqkI2T+zPFe4CEusiyL8IRDuPBANoSbf4Bu2Hx7OxjY3lwGUEVC8CbAp
yGG/cELEFgc3cdTMLiwpY1bMJ57Yy396j496do/WrYQ9hH3NGMvsXlqfS7JJyfQVYqMBVaPgvbfL
0kJ05VBF9VqgqaucY/27kY0fHLujSBMiO9b3/NQq6Eu/BbHG8ClFy2q0jDfhjifgffGvLN5W9H5y
tw+AlmxhiGZwSvTWEGlLJcreQyPVWMT4po2HDvY8E7PZsxTR3Sg88MxXiIpcuVKrJmJ9jJxXNVzX
h3poDYhy8pxlkAo5/Dtvefk6PpiaGW+cEZmQfmzSu94xa12k0IYEiWNc3XNHIy/7dYhry28sX02d
eh+iVEL2mGrhlHHYRHrF8UXAbvIqY24/5NSw/V7wleQmTn3Fi2DXTRWcQcxYxw9tH2BalB2oXKZu
n+T3l+xlDi+L5Dbk3V4dirKTrKPKm9WzOTmEYgDA0v7orBh1nXvjZODpT/ShHua/86YNL8HUFrEs
R3ksNWMdXByYyati/IJQdolXSP1lxfuOFiEJDxnYdHTLJ4SB4jBGzfdvdtS9AoFI4t/Yyq6b2YpP
IUzFcYlYyxQ+VlJ2ithllhIbQFZ9P96ZvS4YH0e7/wj/jSeuZJX653+dltE+OoVvi8n0eAXFYkus
cXKpqKlkZJxlB5JZuuUWoB4anTGU97haghDGNg9qLBaiE0zEbpwxtpnNmLpvOk3exs5EW6j7koTI
TGC/yHrDxli4S+sXwMS3NRKYMQqjmfmq34bGn1+ksQ2DQQ0O3KJx1s8v0Ax8iBtgGRA5/2jsNcj3
eO1IkaDFFtGQ/1QfQBa01gpkTAXPJgRQQCuSRPyRHD1fiFfA2jT3XquIcYoHUFPd3BWriAcpFkwk
PqyEbZmez+/y1jb64iQ6C6vWPK7gsvB9TpzlqTrhpQcxKb16S3wLVmNAcXLKcunfPCb6d2FDyLTD
k9sdV0YkyZgem4t27cHvgJkYX3+j6Oqcl47Q++x/D+pEhX5Cd7x9DxrDJoh3xpd5867Q5twoIno6
HTq2X4xCeLRdqbk90s8aaZ7dIZgjWQ4ocFlgo6NLGc2DheE58wrdydPmhz5PKjoYNmBpN7vZsIsz
IL+SBu0zC4sRoWda2E4xuJuTF9/JKip9KugAbpxwDym7WUTvo8r695SG8JLC+TOXukYaYtIX75nv
WjldxTJShwOmrORH6KBH0sCggUBxd0sT1pRcB1jFD9id6vXO6oQi0AAZhdlXKGN0B7Fp+9uU+tuz
qfFAJZ8HLOZvFhn9UGxyoIJD9KODd1AG6V+T6EF4kYb5NE1PtVyowKG8gpuzLX5wpA/X85+NQ9qU
2eb6E3/Fez1DRh7WET9mKLNN3EYRNyAbrFJxXA4ePuI1zdatCtw9iFMJTFqevJ1vFacCOIyxks/Z
BdIGdf2f3JPIieMClI00J6zQncFc5ILG8FB10EZHpI2vfNRTpbmXSAqtKUL756iBZG3A42GgQOlA
ZOCnRVcxU1zjJWFRTquIBofwb77W7vaUfMJw3QkYfVziTv7hLVZGnj6T4pTxt6SCTkFyDp2dUdiA
oh7VwRG3gVK7mTNPnUQLZPgrb9wzMOHmfGbagI1p1N3n+AaXiOKym4G/QZ9DRPnMtsRjM4OzaUAW
w+wRwUFrhhgxh58+hvH4zrms1YAhG7PVmx53JD8YJfzJGqQA5Efk0Cr8u2rvbENZHgQGjJ5EzHMO
jqvvpzViyuWmSaNwBQgEuv4M5+7UK55Vd6Z3ZRnX0lcA9buHJvlScADf6puv73wlBt6ttNALD4ls
SOOlbmXK6oXzKPjVyI5NWR1Rfe3GhgwO5Db3ouhDjhLS0tCICOe/SIzQ6Jq4YhptNfFGucbq65x6
URY3j/4Dckje8kV/glciS1hfaEBu7mwWdy2ZraxWL1puFJS+zRe+ZXTGii/MSEbpoSazGMbl2wfN
OD6wJTarhldeilPGr4/U+gevYPNbdyInKW4SMcf6En+t9+OeYpXQzoFcuMcUx0nuemqSqEgQrYQE
jKNP9vrdvKkh7/wEzZtf988mz0HFxFNO3T30No4AM7mc7Nw8+aBk/AVLINazv16Sy8m2vtHS8Q2m
ANfNTiYgGkViDHAEl4pi+4dwrifZyc2KcTzQAk9UO0c/TZfoeIQfVxt6ZUZ2uMScdCn1zJLXvKKc
ODQ2X6/TZsAy3btz9d0+wgZx4ak4kydXjEHKvjKmFJ1mm79cCJ2hnAASzHyXlporZ/jQRG0i7nJk
GlMo2M/Lw3eFpKr7nsJkndKWyEBF6Q76lyip+53U9af+vXw8xVgfTp/yyXv9jXMY8F6WMzi/3h2/
EeNfNUleaYgqpbVSgXwfS3KPjoIpjtyQlYbP4Wl7XR+ELq0TD3t/fhSr36pWlS7sTt6aTgtMBNol
dB0vw0E4LEmd610Ikf4yzyKaRkjtpPH1vbtWciHZVBRtEgtxaMT11fcXJxBWENeiQeLUlySfSIMV
gG61oh75wXf3t0MKKL6ysE0oQ0nHBH+Tas2k257E7UMm+O1R3DBWTWpdomK36VgTvlhYnLUMi2A4
ML1oNMMBqu6QYFx+fvmpgrEowbligfVD8f/rxugDsDugImghZNrc6SsL7cP4nOfY4nREeu8ShCOW
o6/74jT7UhgiqFmAN1tjMiKgm8M7jADucSyAJmMdyGSn2CHEDcLzapzeghdv5KjYusWkulNcYf+N
DCjUY4GwqFpC2j3N0kC4ivWX/hpThVcAXNUK7fN1Az+Oofbk179FWukwZiUj/Z9mathHjsuL4yFq
aN5r0Cnnd0b2q9xJsOFuPwh5u7mLfyux2VLC5G9ZWqsRl4DSCSR2VUVxTXBxvGtw9yeovyyQuzaY
5OJ+tg5eQ5aWJo/sENFCv4/F8pkVZMbPrtvaykJ/piEZIdmNNWELp9kffwad3CGpEtKedLTkQlvb
F8C5g6CiNbcmcQeLgh4LzP4n0pXMT+syD9rZnNsxqNf/g3ppiDeaN0o4ERuWM8pXAi8FgDRBQQEE
guwu4T8k77fRNvI8b2yuDIJo2SKFsmJ+WFUIzqYjF0YVDDKqmOIlLj/SlEb/Av60WwuTigWvrfdY
x/kTc+iDdLcZ2sKfXiCI6JaSJgBq5Acr1iCF8WPzEmIsSfF83VroalXP08fc2l4xlEXpZQ77Q9Ty
b4h8zSD/8fCI5BQz1OqMbDGvUTgdJFcO0sYwQnpE8a7a3GBJsqlRw6D8d+AdRKsBw+WYqB1KvQie
eleOVCHLOLLveMa5V1nNOj/mpdqUJvn6dc7ZP2/hEi6MajmBpHGDrgCjcdYovgkFG7ZOYE96KHb/
W5ke9Vj1TRZ8/6wZJH3R63rn7CHtPozGa17s9lNNfxe84fIt8ucQWYu16DHLhtrzT6dA4/6u2jMT
59L0i34AmgZRb5bqqPg1DXMfbmFSFZjSbOiSZEuAnqhaOSRmSw4I5IJJL4989HlWU1og5Iybmqia
oCbrNfZwYYt9Wu7IV2rJpdu3usd5PJP2I/0Av9yeWho/2ftoGDjGgyn6BbddRgN2Af5qwv/GjIj8
1ctW2upG5Ctw8O9HLroKpETXzga4NGkUgxaFGDnh6T4IG+s4pdq3MckBs/rzEyNoyO6X8s2gpu4P
dGB5rSN+kQ7QohuYE3muLoXqAA/7PtxvA3nkSbOaFR+bH5fxFfscP7fyaTbIWEFAuZcsWmyzojSl
FS3vCxut6EnPIBbzNszJTCui7FwyRHrSqHKL+FsjSyjzEQu46k3YCK8LXQREeqmr7EDLYw2zxgtr
3HEoEt0ufCa0sHwRKeL5J7+Q/T43arinKrw8NRSOjbwDCvL17dlb724tMpa8LstdiJ4jzof52Fvr
jVAXRLYyO+n6PckyBwIx5MPsUmGGtbLGWLe0sIMu48J9NWabAIaC9FOo2glFPCscL+1jgeYEdhvA
esJ6x69CrjsSoIgHJhYr1Z6Id9vQrfRBCkk9lb9TSG1HpqMlGv1jby4PkWE33JBljLBO9++qJahg
kkxQcnrUxJwbHGWMswCqlRFvNBU/nAUKFMjhWS7lfW72ITomJQhxTfhfWqnbNC80VF0ViXKDb1Mw
Rl/8DdyQVeHCbRQ2ZoKEW2Uov/uRpsuO5W0l8YYj9HZF2wo/WnqfL8J6/xnivD1GXSuJzYlFRcA4
F+MuWGqVX1jWbmEB6M8erUSYq4jQ4XPiOG7HScn1gquZT79ml3FtP+3Xa2p56a59Pv+SsEf/wWZP
nq/b4R+bxB6z4Wn37cGdDCrKXpKeAPH1xNmat6WClnEa5+WyAJcmuByDlZRct/5+S2Sq7khZAMGc
eCip5LwfFwKV0hOAHDJSgxVyKZCJaxlobRQG0vvaBegbWuBq2EQxbBejderZee+4HJIsHC3TOp8n
bfua0kADeaSUDp7q/jUVQt8Qy//Mkp7TPug/GGwYvq7qU2lXElY/hfwj5OFNR0T9nvP0z7xzKLh1
B3waggcJuE9I3C3Vm4qd6nu6lHMBdpxozRnnUHdIlpM5oChGNaMnAp6WNno3GaosJ/jYLbWOPo7L
Di9oiZsxwP99u3cKMDs2Iqd9eC2/ZOsETBx7SYZ1QKyXXrUcLWJ0f71kG+3lIOni9zPX8RX/IUw1
NTHE4sXv7+PEW+h9xvu2EeOIMJmF3e1ZpZI/Cbsrwt27zkVyK0jPcuwAgkAjSCBaC8E93HxGrqu9
IvTKlMTC7SL9ihx0SFzvdThtoEovjpw4DibbEH79m0IPQIWwGWP55x+t1UBOBXpA9H2KyD+l5n6R
r6BjM44DzkuSmh2vaoyk41xgR/Hxj9Mz6DQxAziLGmbiDhjmvQ5C2kUTIQxmWsJR/sGS64oZTiPX
P8uEVEUfFPL4CcAnYkdw8HM82TtRLxJCI+htolc8nWQURLHRjStYjPIMnwKITss02bi5X4IyE1gx
R11jkNcYn8WqcRi63GffAwzE7J6q26lVjdoZN1HsCdolhJPk9qil2vegoAgevIBVL2k1ycs4cJ1w
z1Sqa7lK+35VT/HyVqJaBu+Gy9VeRHQk0TP/OzL89UtKWwvMWywiYYjsjTwJiirOXpC9qzfpi5kx
QLryJ5v7nPUc94IIN8nH4B/VEpNdcm3GYjDbXGQPmhmrsiYf7unLupOkwkZzrR5+U5gzr/4Y1DHu
IKad7/r1TYesM9wUSvDMwOK7i5Rz7GL4Cs6nzpXZx18pBfTSCprPqSdQSakNSgWk8l+8e3Ym+3Fz
cUmMXNTvbpNpYVQSZvkFGCaJrOza/EUPSSZdMS/pjEaGd5TcilRFxcFqCYK2t+tAg7DWblxoBGLZ
gaJcvYqs/YGtyTnPWJY9FwzQPyGDEqdMJlS+xqXTn89eYmLNyYLPEMVSsG3GTFHJRd4IVjRWJj+V
U+2QKdpO+30KZhjVXtujCbqTuxQXlx0M6XNFQ9s3uc+NkexEK7p/Xk/7iMNtjkMYj8R9L76jNjcq
x2PzzHf7ke9e0LlS7hZLyo3qjLfo3FteTiZYthYYtTdlWkA+9zIfRYe6OF9iphEg/pIrBymGqi+Z
10KBIs7+0HYEhlv2SiMcaV1k2qN7y7031KpF4vL7AtMKrM6xPBovWWDhjmh2NQZTM+BWXR2vXejI
c+Xtbv9WRYgdtfSyeLnFRYir5yFp6D0dTpgy6XOQQNOpFODfbDLYFtyTdUjoS8NcMGI+d8r8LOgS
eGGGgSxIuMcI3dkLVl8sR67fIuMV70XwtKhQj1JgVS309H35biAc++flYiJamH21avb/ULO8s49C
vHsT44XQHTtm2jHRs+VjstkizotQXq8RESDZZufgZDde0Zvr0LkuFBCentRwpA7740PRuv/D51Pf
RUc3+hXSDwbs9LmmDShKvu5AKCkkwGZRzP57srp0hGohYKHSa6jGCT0RCsrazKxPCCLLs3ZDHqLJ
cimwv+iaYlYrVNuOr0PHnsh3S8tTB/QtTiEcBF8LCSCZBiy9ocUaipdRvWslGOIK1Dqa0SqrT9rR
EP3kYrpkG2Eoi6pA+aTkHg9Srv3frD44U6Zy5fIpCW50yNUO27tFHQGaEgK8zm9C5HlV0aUYswb7
H83uIeDWC6cPbgpz1udEPXpTpF/V57A4Kz+ADHPzLK+zngRqDapmDVK6h7I6e9uRXpVscBizYwZe
GG6Xnd6JU8Iok/CAPWYo4XjJrvmcaSjQe4ywVPZpxYk+D3xj/zu1kOWn5G7Sb0ox0VJofVCgUKaU
zaYth8sETh71aaI9mRaPMcZC86QWTn/fccb4O2V/w5Xa2a8NjPUzF8JIMiPqih7Wt3BGL6Z+u0W3
SRisBV39hKk4R4z2U+zcxNaNPmECf8Yf/r4y1K5wEIUFGQkMI3xkC+ACVTQonYGjuo4mOiCTqfDf
fm1CHSJyViVNIomHyk0ARPZApT0pXflXmen+Xi1NZa1j7IDpeWjoVXkiSziiPSq8nEq+OwqR4SJB
EUqbl56QRnXAB67E/72Qm4rOW3t6dXsGAyobsgnlmgWpMUS4F29cs/pYjM7wMaVZVluPDZy3U+dy
GGskGDjBqn62vykf9EWP5ImsLgm60GcchxpvHOsgFzk85q5G9fYUQ75K9BFzGTLQ3N9Wx6NW3GoJ
q4Gj9eujJ9uu/IzgGncv+QCOpVFpSh/aoCWFpOtYennyH2ZPqQ9Z79R5doRkFhslKPEGO5xwQlRS
+GqDFuWDzZR1x8mafvjMj/Rz4DIzcH36moVyT1yUfDsGiumRJzXqPD89F6PlQVF4qUxbYgocgpOH
G70hmKh62YHnGRmYCAhM+X5n1BpzSgvMRkH0J7V8/JIJ7WFhjxsyCX42vVMT1+9YBtq7Cqovbe+X
pM/DkVLp/T09GENYtuFtC8d/JvPUWAsD/7ogSr+aAfJKHv7fixi+z4qWzGI0nO5EOSeq7HIr0TcU
Nousm9hPycEfzc+Ml9j1ZGyuYiHjvgmgamwRH4NxK2rxQjyhVmnoAuYqQUbVEnSjR3p2ai1oPshg
nnhC44tsEUXAAm6jhIZJpI0bcoZdXt2LGQrzcYZS6Kv+/I/Wzx3KnJ0shdab7T9XGTseA5dO85LZ
p5qPjY4aErzjnH54Q+/KebyaOZUWyhiuVin6vn5HdcibzvOD/ZLRMu659y05ZibEzLzt1GAuMwc1
OD580rUbBgREYJmD3n6e6JoqEuGfT5y4A7yv4YKEEfZRTW/RPVXIM+fOwrVgjooFeXREnO2oZalY
owB+CqoDAPE22L1Qm0FWI+/sJYuHEHZINW9ozHluMSu/iSovcVqcgT22WXOkh/15TYxVp93WB54d
WVLf6Itc3hFzsdtx6Nmle16wpB72erNNFFxaBSexKxG+ur9XKyV24+Nwv1gQui9IY0Gb4NRlV6k1
bDicfUt5ZXwuCzRk/BAHYWms2lh0RT3riijkh54RrqLRDayy3oGa3kNn9LiHFWFoARYMV+DlQnML
3yVIvFxJpKqeUTHEDvAycP7vZj9IR9M4ypZI78ZYzhHz5lhA7dJWKocU0hf3j/XphqmTNsG1CsXq
iRr96JpsHuuwuXG+bDLT3EMvFthmNB9jBynP3HPEmTynfWUJBRkQ503AdUikp0B1Cr0M+pJLAYxZ
S/JZ3P7gWq5oDVpHByCenYBeI9jqa8ozHW+n1HD50px4dD7MyYHlfpApbVBLQf/sduLzisxZNVnm
g7rMqToOLIbbNtud7082LyfFKzbLq1NjU1c6c3O409JaSS6zFvvSafev4ZYzW430DnAQe9KzWlun
Jmbkjt9eEFFDkL3f5J5raOt61SXjMTHKnJi/SMPumgzI443EmLA0bUkqtd7FnVLdo5eUtl5GbmCr
/xTxE9/u9t4MEKl452ba7lj/kZXHuap1Eb0QA+BF0HJ9JkJA/ezMnUZw0KCrUKKAUZqOixOZ3ky1
duUDmx1Taf5lS9gO3CxoV4HufxJWSRAGDnT8let9zLxDCs/akuu/Fh0OD4+B/TNZlJqZ53eMjHwC
ykN8cY4meP51KcpQHf5HSijTlpXaokZ9ff2xJ/C5VtY2mbvfYw/PuM526ohXSMGWVcHhqTHzIY4P
DGrLH95MDNJyNpq1F0peMxtdHWUYAErizZNlC2OJlbyWV9eDCfjcwA2MvCUobFlTtLxp3xJO3LPy
ZAQFcMWplV67kA5GzayE/4gi9gQm+zjOvrk7bJDPq0WIdnLelDAgptzK+UQiwCVCuqHY580Tu011
REGxvlgcPJfTP0jteFx5MKCyEKUIZS3Tk45WAdCYjoFDv3HYLqkcZjLm/ZntZc4L1ReenRIHI3J7
sGC3plNf4iqw0I2LSKQUubSeTN8qhnv2+OSjcT726Z/a3fPXGdbTMBgbwqZWcODXKD/4MfSRvStJ
ZIZF7aeBq3J5SnGT9MEWJ8J1tiRhOQ4AmR0V19b6kE7xJyV67IHDepqUjLhfzjKX7v4m+CX4fnsL
Ck/2XU1rk1y7XMMT1LteVtkqOUmNeqSs8Gtxi3VPLmwBTZxTRLM1a/HidXOS48jWVHuVHaJZGp8w
PrAA2KDytsGgJMr37qe/fhS+sep/6ng34/JtvTbbAPD0pWJzJSS0uu2bP3uVhHczgEvYGzQN70FI
GO42Drca5LzSluS8jfCW/9LJimaMnqZDGs525hIE//xLn7F7LcK0Q9gm7R33Th80HrLizggSGKFK
GnzNGk+jImghOPjHcOa5qszubnb0wCNNLGTBRXDcodfk4TWxAIq5Y55yDt+lfIBEWYnfbz1E9grG
G0adAnCZI3FmQGUSsGv7YiZHksB6Q6CcoUwCVGN3/B+mEnpH8uzCCgnSJEHzRGk7fdQDbO6ba9Yu
2TJD94fLO/JxENIXRyKBRR3tpRX9PCKuRP02sZxfgVv+DfMmOKKpz3ZRwtPsGWgV5wQdQWLw+LRs
MTRfge81RNOePbtbj7YmNsqOK5r3n22ETn3KCioob004jn5EkSjHF3T9ev+VSrTl79MdgxiBsAab
zcuKx6RkbT6cR1OHfLIeX6tLJZpovWYyYvxqUFrWha+uGrBHemiKI9WKxskRuSr6H/wFBRAzZPG8
r7s+uJcIo/TsYq5RmdWfjgjVwjRjMDLOvBX4Mg4xii3zCsG4G1cSLhpwCcUm8PUgn7pZe9YMa3Hi
A5Y6p09DCVtSeqP6HNCX6qgrx3wAxl9DcWtH2FQgV8GN/Bddb2IuouTPLsZZ2yaneKf4S2U15EOQ
m+Mq0RGpG5Y4uMJS1C/hbFmbRAXLurlyjFgUE41m5ydlNYBRKMQpD87kzx6TbykzaYYQl9pKcmLW
NFrZoI0wJLNbc1ma2pMxBcXdCpY9Z60s++yugEwjv5MpPrlgY75PsSwoo1809j+Dl842rtUQgQ18
qB4WvcRDRoyXsKW0s+LI+UH1KkG3WpdyOMy0oXX0KTzuX5cyKEsBXn7I/pbGfNrNtRUohkAWDkr8
19YSiCy8gS5HMjx2PoKMFOBVx0grsO4khCS0zJEKnM0lwC0/v9t7M7fFCT5J/z4hf9V61sUML/jX
RACtY9wq9piVbMoIfrhNn5gJnz6/s3NYs0KOtvr9JOIftuPCEl3yRj8N9kOMhMCx1F2S6nuala6t
G/aygKNIuOXtjB3qkK5BInhx/ORb2ilmxoiAUTeofo7PGe8j4lFe/9GcnDbs8kWalYpOKC/pNjkj
nPaxgsbB6NHeBLVJjeeVmXjKV95LmKKeIF171tA5N9nKZvBgaE5nAOaAsPHpqqnqNPPFsYk9yAXU
zO2ZGStjFgGGviC3nblQOhHz6FhooZm0r6FvsNqX3xGVvrMcM3Uh0qx3SFgIzgOC/jhpt2g8SOwV
yTM1SwtaCl7v0rPLFySnRNG/CMTnjKz9Nx5gxJ2aDSivDVcQtDW1Po7oNKWRgi798ax2ng5aLGAJ
LAgXJTufhIosLxFmTaPDk9Dpm59lafYKrhImW8m1lDpJ7CDFlEFrW/SW2VqNn4sVlyd22xECaP4P
6kiwEiuM4ywYKxeyuGcJHKhv67XJr7dKM39jFmdQwoMl3hUIJFeayjUxXGhFM3cbdyoxF0m1Lj0Z
L/O3qQ66HR9o1MMb6LuL2wXGBTumYAydkH4qlWim/VhdnixmWQkPOJ5Nq83kLLw5WovX34P/NCsN
pQWq6NAvNqJX9NMjfDSZsngx0oVFNnEwvIy7JTsGc9+yvhlpbeSKsfNy3dPuhDRSkaLtfzsxsWYs
PclEX0Sd7+JvNJ+a3X2C5UYprHRhdimbY3ze379BAGE0ZYk1eULZgwxY8a/vO1r1DvFgjpM8FCeU
C2btvxNckEsCdKmfbzJ9GQhgPbQTlP/MmWucsNtG321TmWGzhTPVcBG9bQ52aRKGqWeefyFzFc4W
HRkFCFAxBHEt5P49xnJ8UXpLvfNOYthVC5/anCs2ot6PVAkKt9cNtrOHmfzsTJ0wNvRe+/P2jv93
2BJpYKj6TjT7Omsagp3U3r2A/tM3HjQJylzMSQdoxZ38d2ijEsvWx4dElBC3Qd0RnU17MYv187CT
FuYnh9KneZreZwC8x/Y8xSHPI32ZL3NZ9ohKWR+QoZHTcF6Y+x0qpJojXy5M5a9vkfq5APMRqAOG
9LBktXJj0ZQQKuyPYg/yG2EfEQKQ9rIVetIfx+DirFjp0M0IA2wHi/IYZvCce3m2oLqXSx9973Xl
rwMuemF8UKTYr9+eO5SBnnIhzHK3G8LpBMGm8AbqTObt9Fv9e1rwFv6m+tO3EH4PQFcgDr8SYqBb
8odJDDIE8r2rs1FecJgHH7QJlQk3tqTGLN0x8+JXerMdgBqaXvdQOOpoverRb4ynaMheZBnIYr66
nkvAbHSC4HdRbGJ3glar8JiPNCg7sZL9hh/+txYfJbKB2Bz23yHxZ2BlDc7g0+xWQyZYufUBRodZ
1OCpz5ss/gIECZBkxjEi7dLp1iAdaSl2zIMWWkTJSLXZ3KmDmU154g8D4nI1FsOa0jnPkrOj0uDL
ihJxaRXDUzgPtP8UQOFbKvng+R11+I5A2VyeA/5mMOY5W+pvUAkQlADaz4Hk0lV3Cr2InUo/AbbC
VHzfj5HDLUtW2OcbiY0fQq92uiu8kNXUsZRH7sQ76Yn/IDqkmaHEKSbgXuDh6c3kBoh8SDTCLeUA
EZ1QWpVVVI4Rm6uS1QhVWeuWYWcvc68LMIAFFLsEh54mlnODuT6vKBBlCYybjlP8B3A9AFa9yzdr
20W9rhGXK83JFu2vnP78nfh8Baz+izfs3NJJhJj+0SKviGqalAaiYdJ1hW6KkBSLw+36sxNBeL/d
Vh2CWgH/+rLqqNSEZAAZOed7loiWIN6/i71NgqY8HVEJFnsXA+rand5kxX1TVBOkOH4sKGfNfCfr
Qjml0KabFHYwp7AV0ZI7PNi2pXygFBzMioVEDvxD0xuktzLkS2/TsVfGmHb9igLfuHBdJRGxPTwI
YIAYl8TQJDLneXvGXITzTUchF3yNxkVEGX930SHfuIHzxzUv9eYO0xNaEL3DPapz0xqlXEVdc5gu
y5oL6RpKmfsC88lD595J6gZg7Zr0nxSz7eCHbPbz+vkNRXxGHPq3+/cvnqfpQao9UxIAUL8fNGx0
DqAz/AIwkn9+5rwrVmFtsIML34rsUCtIbdWeon10XuhfpbatJd8FSPm4rGeL3I4MtA3CmSCbhQqz
PREjwmxpdaMgtT0RCnFaVpbDQo+snV7ALdAGo7fXz0JqEizWVySsnRVwAGQWplWHbCv8c3uWin1n
FLQq41M6qeYByz/luxkmIarRbmflITO0olCePKq1hcDKVI5wsAdXgd1O6w+XbCPzDJhoJIslI+Lu
ktkuLTH0GtUp6mdRBGxr8pU1q4dW4x6o2N8CcscYpMYUmOkV3QJ8A6zfyTUC//OubIILh9D3y8eT
XwxQJvOo0O+BFRrup45ahytKZUONl8cluQE/+1iWNlZbE6AMY/vxy9NcQBs3ruGSNeYxHJURpRAb
NzF0MCfZYLKwqyIg4cj5ELybnFqg2mZlHwUm6s7DC++ZuOtRD0f8NiUhqy21Sm6JWsG1fbQ155cf
uBMNEXo6XS0XyzqbUkfkb0O7M1T9P7EOiDZfnOfWZnqA755ljOo51Q02t3woj2J2+fQ79d2LKCOX
+kDFHRRRB9mjD22euHCg6Ams88kr+X/pOYxhyoJ/rxN+/byucJLu0Wxu2oWHSka3yanRxfBYHjf9
geJy25BNXOB41aXZxkf5EPJOs//qwVvkF3DvWvSGbH0+rYIa/sMF/hVwFFor/iFOZl7RqDDEQQ8j
Imc3SgcVVx0SYsgOiKqORrAFm/UKUT77ZuLfg7NM5dQl8xjp1TNXaxhxIgRE+HXQwvpADtXmyMC7
w6O+clgaNekb6k8El0Yx0YTlFpMeCZSjvClo/e7ukakP5tJwtdEKT6jgPEr1rzz/yHytHQiSOTBV
XLbMu3mIuELc6ChmbXwmFgCRHoj4o3J5eUVbbu9bE7anl8izYVupN8c5yTr4ftEjkt278egrzNYF
C2FYWoMB3y3MgYg+LlDSo3vuEjg9xF3fVqcIvmrrOZXLojLwV0+vqlLKxEbre3xa7l4IUNgx0wfB
brxfh5S250as21gacgW7s1j+Z7W7IzJv+iNCfdAFTaBp0IZya66hCA/XHt/rT4PSndLJPsqqPWTL
FnIKLVgdG/lvzq0C9vXQoaF10OerkBkYwYoNL7y8ip9jRIf28zuu61o29YAObdET5ScpsQ1Eh78n
WkkuVFjWWMp96gXC5JLLdQm0NuSpmUMfHO9ksMsdr7Zb18rjpl9FhIZNlNjCimv8gCmRaHu43dT9
oih+BRLFd7lXbpz/tLR0DInvks/U+zlqEKwQlvrxsWa7qF5xwSXePVaa0RDGVqIjusnOW2ykJyHg
ritcqmz3ALL4hrmQTri3lt5J3Y9L3T2TPjZct5pkD2nZmZKRY4rw8PG7yR3e3oesOsyDP2q899DD
rcOjVQbl1ZRbAU3hVqchayK2AzJntq22arNwXSuJV8JoDUdhT6m3d97xvOfwB5FvfbldGDpQbErA
Q075G2NUI7NE7PkBNWmAh5HU7xjJa0UhAT9X54LSfJ0dKRVSFtwikOk2DV4XOy81CqLnh1jDoflc
+mMu8VuBGxTDYM8dQy8CsLpGh7ILlDF785OwPcb4HoK2rSX5waGi6RgRBtlRwTGewf8BbEJnQEIL
DCvpawMDiLixWEdodXiV5Q/SEAN938s45fSFkqHdEWU/n1eryHAbH5/ljCh/5FAJKuG0zuc/mZpB
DcuHQ0Y6XMZSPB3FmZ1wf53ukuG4E+CYZRh5FtMJ/p1Udv2btyoxzbjTFRPYxT6Ecztx7UWg4Uf0
iOVRj9bwBelpG34cpKufhh07qc57P2HK9iNgIy2scZC+C2fYIlc27dYuTKtigRMSHqXJ07RGQT4n
DKTVOsYc8RJ2Z8GHSKfeb5F3VgD5H+NlnBy61jW/Xeto7LXrKKFHW1LHJrk+7BJ0FMafRkgqC53k
e54Wc/0LhrKqo5uRIi5E/XmBi/7OdnVH3+/3h1YWUMLdTlI4bz0KU9HCfODGeYT3FZSYgQH57Ht9
dv1sXHRKi3rjSTy+VFWn5OX55JTMbzI+ZlnHn5+gZ5S/5IE9dttnnO6cVDcJ5eSxKSbfzbnw/u/2
6NbayAMSppfZ97yoIW5TToVZIzVHx7niu2mybkVd06TFa1ddDPt6UHV4S6bpjgZcuJJc9Uaoagmy
V5NbHO6aUwRdQCbwTSdZi7uXRCRnV5sDQ378yJHKIjGzvYmFvGjR+4Ru4zAqLQ+EA9tudajNdE8V
iOelRX4BryH3resVJGl/uIGLuaPkhAJfK+Ot+BsjywZd19k+nFnoQRc0coA/Lzh7BcaHN/a/+x9h
aCjTJrYEqTZdQzmKk15JLVxi7SgJncRUKxbUhsDpJZijQA59Rt1FXwor7azGDeDRm1H2/+z8cEru
vRCa+ly/ZUo5hhnO2wG/CrvFF0zn6962XN3LhQrHDn4Q4FUbawgu9njbrWGEm2VxyiG/sqcwU+f+
0dxi7EKhiGntoT08rwW1LudTUu57fVLDuj3fA6iqPJUqsTEGFdyXIey1i3X0Aqm68kH4dDrCu+PW
5GJp21bWiGh7Po6Wz7McxTt/4AuCqx0F8cHF6n3pWHcZ7UfacejaZ2GTX+Qj8U5tJHyHizWol4Hf
7+fTLLrEqq40T09TxlQ5Iwr+TR+AtcZ4L+VkON7J0M7u0cOQV3MXwWawN1ns52QrtZShtCkZiGh/
dT6kfg30VivzEIno4hkfcA3jTFW2T1cdl5VK+GIkXrTwm7Cxg16ccCJST6D1nuPS8ndSv0cesO0Z
IQ0hJbbKKdR+yjSBSD4OVPOce36M9pwNHEcYNdzaooHYg+P5ZTWf+uUT2fidCFpfW27Q4Y1bzZxz
+QBkJgehKrll2wP9hagxkOLKK6NTRlXF/oSeHngFxztGRdsLSQRzkTJiD4ygviiF7vrRssztbrm+
0cR/lusHPjDMhwria0EUYHZ31BHdzFHxGxuLG/V5RhaxckXeenaKW2uw29UQmtQntxIvQLSxdEKw
eh5wS8sxqqiBcKiluDuur4A7lx1edGpqIQ4dIwQigKO+XABwULA2AfqCLud6Y6ny9VohVAXBOKcr
4CWKbe6L/9jhrHmO2GTg1lU0t+sYPRblbAsRZrtn2i85ICZfRe/69KLmsKycq4bl1SmZIbYRhshp
SCT1xSVRfTKPgR7YKg2zkwGzgpJawU9e12gJtasEUgS2PYC7JmN04dFCfDjNErkTW3uEOb5GKlc7
d3DNgJUT9N1bcLFSCOQaRpnz2PFrlN9tbgkLTORC2bjiYbK/GgGsPogRjXwBSX7NlRj9ER3qj/16
n9URAqF9/Ffzd4mhoLdCkJnQZJ+bEeoDz8d3tfpRSAZeI+rPZkcYBgHiFZ1uVfayz0vR1IZU23U/
UyU0rIvnUpLKBRYOXKe9qZYfAdoz6u8SnIU24UzuPuMvgAg7YjyNNxGMSuDAqqH6zh5BjUZD/Nve
q1TqxwbJxshi1VsR59KDlA0gpM9c1VSYw9HifcZB4WqBL0BRLLCO8Znvs1lqun8F3s85I6phCwV2
wvcfZfJTmJ6FZbmBm+DRPhTk6b6DlyvY38XpxB1jrY1DjFB5C4M8loZYL6yueXJAT39eMmMpJg69
v2qHv9WNf2wn1KL5SnhiGEHj7Q5o1rcAaNSg7AAdHZGiyW0QVe1YDesmX3floVDZNsV2x2uoRjCu
E584YiUlAS2V4gDsVp0ne5rTe0y2ohE8wwkQWOFElLpa71zw0RrPJENmJvLnMV9/LfhGJ0jiWuqF
qCChzKy6Yhjdlah5VqVoPIjnwSINgKBbMXxJbJ6lK8MOuf0/toAmWalnW8kTkGQu+k2Otn8+mij7
3qMM1fLZ2Ir7XALcWv0vyOQ9x8Thmm67txesfDD/Vjk5im3blFXzDNVFiPtFImEzlvJSUnp5t5fb
rdOtThUBJKlFthfnVG4UkHpSr5XQCein/OMtqNs80AOrP4kaRsr6TvshHh/dyFmnbyrXRW138PZ1
v2M0qtu4M0lnlbSNajvyxlSHv1TJSCXtptoFTCFZPBbicrpuE5LqwzYVUbhYL/Vi0/pPfDVe9Q2u
El6KfYTDmZSs57oLsQXUSSxO3ll0wqPT92SbfavLaCq4i2rQvb3KwMntdfZ/FIW2uwUBWxHBkjps
0wfHSa1RzPmQGp9/WyGaNjQTVqJcMrKdav7VW6cClgbyLu10AkgoMbBmzWKoMaU6MN8P/FnH5Buj
vvGfx47FNqu4tBY7IuE832b4OBLr7dKCypKo92AzFtZY+jZr5hBqbyKPi1BgF2nkcDm4DZ4puUzT
aaj7zBls1lC8CJeQTTYX6DawXLR1gOHqMX1L5jhnCLG4tX8BiSjPS12iUNhaUwQMRFxjytsGNE3a
7xxXJ6bWWuPTXZ0qXvTTJDl8BoEAKbRrD60o/Du8KK7z77v5lwqH0FUsphk62k6XbzX80QP0p4gG
VaJNnF+cOMhpF6jpG8FemZ0LhOcexbSmcJkQ0EciosBHJYYg3usSAtZ01RBWVd18CBNoizZzINeI
Ml2FT/Y0rYcokunlwmZX9pLXDpIwlBMOimcTVf3BFW/z4Yi+D+0+l4gwyGHgpm2jqfZYRkbiY7t6
sQunMhaH34XliU2Gf0Po0xjXsnSD0ybiVKUlUEjaz63xURozVOLW/8HME5N4z+v9Y8W82fGMamO0
PAFSvzECfkmNGj7P+u11ttrWMc/U3NdtsE2JbGp6f6sWUUWA+KMgmcf/eF2dbuz/60v9qmJNyaxw
uFkdZF2a0D7Xs+TxcSxv1LOo/xsQ5U66DEZyhxoZBjkz7AQLu45kDjVjUCjSglruzKwSO3cRKWBw
p16scNE2Q2NqstIfT6DUCZ24NIyUHUJF3Ed5V39nKfLlKTgyMdoDDV4G1WscmWS80s/qqLXdB2MQ
3mbkA5xESVSkU7aUspToC9oWAiL9uHneRU2/F/30Qd+pOk85dFplMcxiIl5HiS5xe+lTO8OEsMlI
BLZ0UFVdDXiksXXb39OcobCIbyjN/ECbWkNxG1rQqcplayfBfK34r9MTyG+jzK1Lm7qlKg0WAARx
QQFZrFIjrThrPBNz+MDkQXiB/5RjjcMr3NENdxQSOhU56w/P7F2e+NHEbzl0cK3ug1qIxXJo5Yu5
joqZZ5EEqz+kVJ/letvF3tGCz73RsowC3+9zHzKrPbojEc4tXf1sE5dk+oJ9T/ZwKqJN1o05Omtt
LLa1NB1FAWdXZC/3lqH4WN7DGw7rF/KEs5wynqCJxw5l59yvBZzgKR7RuZipMmxbO09tCfrEb2sI
NN2Dz4ZuVTs/V2FCYQl16Z2DQaE+z00X+6COtRKeuZQoPUJ1FgQDJGu9ZJ2h1k3ogk4wJyx4xJk9
iNNpjMSSl5oUxhRy2VdS1t1rCjirepVG/yiwr1LTz08jqdegQhHs6pspx7KRcB3eGACES/yV4yrE
Rd1bslxsFjojvZvPWXBWNYFyQahtAKy7woTWb/XISARFyhoPlgyqcFsJHaTlvseqpNgWXBXQle5I
gehd0PZHBa53uqAmuLUBbqXa89s/X3WRgEYYnYpziY8lsCEQzdqhxVEm0+8iPlKPxkigUCSDaZOi
87STFWSh/t+Due3KlxkK/q+e0AgaXZeMfODNSz+u+6fVPU0aG0Xn63Kjy3ecckcQidB0x9RPpHaZ
Gz1vPTzCL39dEOlfFTmcLVNgFhThokfF+OBOM3gQdS4EKKLXZ20+uGXaI42hoBKK22G1SJ9lTpKP
wPKFD2yQzAX6n1E5+CMs2ZE4zblbadKD6Z1OAnLfRq23M5zMoqqi0qe2BmSk/AQ4/Qc6yUxsKuAt
4HUVGBuNM17265hMAenpY3+1NiOLidPADWb6rh9Rm/HqFIAN/ooTsGR+GRHdlEhDLkHtE5MVLtnw
E5QOlT6g9Cth/Cwzg308nW/bq1bj+7cEwpoUqPsqNtCMiBCT9j8iPsqnf7kaqn5M86aPTmQZnxPO
skdAMhPqKRgsr72mymQ9Bhc11ODJKPr2zA5FAbfl0z3ZSbATaf17+hY+vOEtpIe1wU09PlaOlVgO
cxnj5vsporyb+20B3S3Z3fWShLbH4N3hbVbYvUSZr9HxAmqXnadWGZBgi1iXQRU6/gL9ZGxl4HZk
M603M5bioF5IG+h8rHDmZm8+wkAfEK+sVGzJo0pQuHa62QuN/nDHKl0WSqAZZ2DBaSUBfSxoW1cO
bH9hyGnEb4ysKWXmoCQwnQWEaxlyioqfa81J1cyIqZucGGfUUKQLWxyImRgQpi8unORiUlv516Rt
O1O1Mo4VtnsaTe1FGQpkLG9RjmEJ7iJ09xHIcjOO8RZDGyKW1+Zd0xKZ4cZoji+uiXm9ktGrIgJ7
paGEWT390wm5cF1WUpNmiMgwioCll3ZPJi23UbPWVS52/2s+x4kqY2EykFSnw87KPwG6yWSBsdX/
bFzsEh5LgZZb0sFP/PhQLuhgg88X9gU+H7a5tYbn3pDC9GdwtUSykBnIZ0qtftIvfkMw75pZEsPU
Ks9C3DbhVSzni28IWQ1EPnsSsQylpd/DL4OKFp4Qm/CDtP1oogJaphGmJwYqnD1PUlqEn5yx0Wir
pKQWruFaS9nf5lLddg162uOQxmlN9qsE3NN6ZgiLdDdmaT+mUUnKuAEuRSXIHqc8yBI5He0TLS9c
ZJL0iJhPwXAzvK66ZuUuYX477PoBi/WuJbyK0WO6MgiEqjhRok9k4eeKdJraILJcJ11mwlEjO36B
DjaVs9qFzSEwZKgDvv4W5TlZgC1I000Tj3BndcU/g3crsqlAIr5MdwcDzAot7rQFZEaH8ZQgotQm
jpXOkjVpDQCuSLaYtTKxVEXP+XH85Nt1cuAXbR0Y0bfbYttYafjZiMMK1Bxm7wOdPn7zfXRRHpxj
UaSF0rbbOw0puaxwI7CU1PE0RgJTObbMTYFAjyZPJaFAQDcm1yYhS09V9BScP5cG11KJ4z7awZS3
FycJ+sJhw5HZ1rOU5hBndg0a/AMLtdWYKEqUPn7ZmtiTqCNoU3zp14/T9dmX1lJovQTAY3PXPbES
awAYGPihcuVYvygdR42UlRDixPN7Az34DcbzSjjkHSYxysfK3e3/EJIlbSqARS4z5H+GqF9weweQ
dlDwD7ih+HCNLJ4KS/X5C7k8NJSKZd4TtnnlortkusYLVU+9UxRUrOsRHiJTDfpUiUbcHh2kxt++
z4x6LwhmXzyQXW0gwqE3Dj1s2EEdp9Jr6GMNdHDhP0svgG5eWOSM3HX2Uq3yj3MPefEQiFHjBc6z
OWAyH6yyi4ZjctGQEtPLV8JCo68Zr3HzCvMlRA4pGPOwPSJ/Hi4A1PswDk+747Eqqk1QPq7IvoVx
qK0DXdNCyTyNFlaM+jYRjVgDlY+jeqhNPH0nqst5NEnbSZDkd20eiB8zeIaugLCM5YQmr/DJ2qEp
xXRuCgoerOgF6vZaOzTFHJ5HYnFnfZMaGDsOB+UbLTW8B3K+1+c+gQyhKZYjwN+hxUgBXpIz4Y0E
oM7KxCnCydtf5vQVX9Dt8lKl246HH/jmLjPapRWbctxBMpZI0r9Q9qMJ07WSKLfgo5bSzGJDPnhr
0pmz+xVAlQM3rcLXcqKJNqW+LmKIukhaGVEGDToMv7s2Dbp0OohBdqhak6Ym7kRK36AuD/0xCNID
elcTe6DWJXapNSetwgTYyU0d+WdqJ62h9fuOldIjXCvpnw7gEwtaHAGmvnbkpqbqABahO6LHh2uo
X8rDb8IayabZncAg+q7GMfKGqKjXV/XC54mmJG1FJnhKv/gNBvwyDVUXn4i3+JWSgYZT1JKcnsNq
b7W/lahjRZkt1JwH2KXR2lQ3oH4auf+NDyGSxcGOMZspYHTze/53O3iiIxtllXzW9qUp/+VxqD93
9vKFh/XU7Vw/HoE/xVOlTw6XeXm3e0dkTVVd24ySziqrkUb00uzF8tPCUr60bASf2QfVpz9oJ94u
aJlIqAzHq7IhnoS1ibgkfZYvsN+wsnrW4FUARb7egq8vCpsPhiy5/Am3JB9YRWnZvENmg+3hIN9p
wMlydBm88wR1VVuV4frHZFQD+z3i3Yn4e6IwoKNQLpDfT2ggda4+ExbKYOjkHlRc2wqfneiDmKbM
5MaMx0H1ManwqEII12nGYxg3v3BzGXECSlPFYiTPy+XlEYjaz0O8IIDV+J5N+5ycdF2yUo1Hz+xp
K1QhKtBip4OMH8gpTbTu+uG1P1JYM6i3EiOBwgHcrwgdfkp7Ulg6xJ8ePVlvac3RSH1lfxnWoqhU
veLTfENXHE9Q36wOy7q1Jy9uFL57OQqqR32SZYceVUerFWHSyV8uZ2KIfviNgGapNjc7Gbmkvj5G
bkDVxsJf9aSi0JpblrhBFTl32fxyIs9aoQHOYyYrI1tmAnbekbhCFtBW2dcqd3zUhieLaCKNrGxI
8ZCeFeVZOO2Fu/OuX4iZwuKP7avzLA++O4Py8bbUcG+7rMxjXUw73FfezcRxjEQUBJeEjI2GT3+d
Rg4/jzLeAcZ4M4hHBYUR6HbRm3jG6JbT+Afez6tgbWALt58DvywFC1Vb+N514lTywfDbN6HSLxFI
D9RfErcNJLMsIAcTSm5qVyJWsUpf3EEDsv/GkhKGSOmNH1r8ARa58qPF0wUdGAbjsXjQR1hfIB/V
5PPKm47S3bypZKgRhE7uRZnMx/BA01kD/EwoR0Ik6TZdS0KEx3fHOuGXQyiPQtoU5RVCj9qm7Q8+
qsqpb2dw4SwTy0LcmmRUKw4gdWfSGT2qyUl67AxSZveqTQxSD9YSSBwEIC/YnSaJRbkWBRBpBOmT
x9OxKy/2QjZXOP9amnzbzWhcnkcrZq2xPjjpEEm7IaSqSoqNAR8rwDTZ4ci8QIey4u3VHJvrVCyZ
lHPw00n2RjlLwZ3bSjipWoXiYCry3ljV8Hj5mEWZ9myXDpAk4llDhOq32ih7jDKR5L6zuPf9/E0B
4gwMYIlPtAqysSm6z8cUv0eFpCJFAaScHPliih6BiJALipOZyRbCDvTzfRK0w4GQmU8SN8Aq3MmO
FDkWpfA2DgwKHmGG7u1SzMPZcthwr2RYwF5HDsk6zNXTDzvHLUb45hEtz2/7slcfAHY4vyDmVPlD
V+njheiv06/njF8jStHwOGaDdIv861x1Y7/yhuI7b4V9iZJgXcQx53F2YaXixa8SdijY05fqkz+y
iTijeyO1CMteRfj89vYTwQCkK5Xcwxo4z/fugRaHQWwlT8/3L7hAKXauNnxR/PXHCCHWr+UeInhL
gF8K/mMZWbdEjrDQ52n80Y/toAI6qU6sF4+BaN7IrdYDNSmDX+3YN5MvS66HjiXwXx1Fckd4fY65
/P1qF1sTIeRUQiBf6VJzmBGl6Zb2kz1leYq/fi1LInOq7ATlC9dqksNcOrezB+9vqJNM354oFk5C
e9EYexLr+a80zu9biYZOsZtqWW5wB+oN13aAAJpzjCTPQ5VxSg2mGQsPuOyN+1BuZboopH4JCc9k
WdCr7NdKeBQrI5nFozAto1gXwDSPHfivQAn4FY17KyBX5Unh976/YmJbqdnKkY8IiP2+z6oXrTF/
Wptjf96eL6mF7h7RwsJOcvcUMkN6oDMSJr0HIT4p9xs3RVe4IDr498fA4GYtAhXWsGJ3ZEF5ALyC
Oupy9xTBVbiAZFhaNd2iSQbxqFgp6ZI3FH5n200ssgBum3qahgde1FkScBJRW6eC3EA+EA4B3USv
fG/JEvsRtSoqvHgoIJHbbJPdH6S2HblS+DE+wjl40jhMkHZOe4KsoXWHUDyHLc6xMBkZBu9GA5er
LowgVwtFLQ/SaKN+OwIlFvdv5l9WautoXZQHwejRCMFCjIiXwpVAvlIA3fQ62xNRyUxoiHR2RlGp
CS9a4nU1ZnuCHYVpY0n3H5HsKck1Xl7yKQrpFkKfs6Qh01HLrrcJ0hxu8cPlENng5WM3eN+JDbI5
PPi2UnrzrZ0DKeXtVu6Ls113ETOX/vq7VZWDjGLTmN65rBUpjZoKh7+2DkZLsFb8UnBkcm2aEKxl
XoezpmnAhSnSYGc+juI/e0G1tbZod8OOzDwFMtRYbFiLUteDvSqZsQ5r9WWR+G/lfFTaMBYI5ABW
V3ooXcpJ36RwWYdhN5FWK/fIsijExcKzEvMKB0WO2QYN9+qA/PxWVwCJhNqLYjWFNqwAMHHbrzHc
6bnrHBFQJoV7MejtDTUgEmPrIT2x47kfoNE0lqYvbOE75xqgFPpevwR34RhoCeCTCCEeZy4yUsn0
lQOzTyxm55MFhFs/lW5YRU4sudC6A8wElQwGYwwhA46ZkTBvDm0Yk0+JNI793ts3qjMeL04DXj+Z
rY5YL6mDK1GOePvYnm2UnD3Fq4+ObDlHVC3oV1H4cLMVxiQjKu7qOXiC+msWu+OvoHJ9gRXWZ/r5
053fbP8FcGRKAmb/MAuf3p/S0/PdNqxphPf0QV0A14X55q/EDUWbHQ3ESfALx11qCILfeg0UYrbB
RliNTO9Ef+lV7uHPkAwqqTnwvH5dEGV7lBE6NvXEX3+9uwP9oT0fiCgUCRbfavRK75bnDhB+wDru
QMmq9ujpnLtD4d2ythjZDpLzNWYyAn/+YRal043fvXUf+aLMAhqYk4bAmRSJWaXjndTsUA/OUzrq
dRmjbiqwkk8STJruUYGttaLGH3kQQW2pmKy0rpzNkeb83GvWIrLjp8ZHXVtuTaKcsRO9DQXa7Vgl
+gmacrB0caACXZJPZ9rvInK5bF2Nm5cPZooMioqU+eQ2EjIVmXZUhaPWJsmosqtUQmnj4LutGTO4
AssAe5eOOLdkzoIUp3pBrIj0OMcZ1XNa6llG8i2/Znhco+uZGewXl2J/ajvlci6gQ2JFl/feg6EX
02OWIuwsUZx3CSOy2BoreXFs4KMA6pni3YTmX0fw+k0rIJFIA1PmGasFhgnVFn5GibPYXPLID+7L
V3/2Z9M+dVR8VeW+/hEMoHLGaxgoYOrf39rcpDbpJMIXcluS6ruYOLNXkBauCqNowadzF0bw6Olt
V0b93KcCd0ofX72XXWNy3Ub4+qnyaPjgZbCUC0M7l/KDc4Jh/X9XA/xA2nr0E2ORvSMR75RiKJUu
FpbPyZluEX/7K/ejLKPJfPntwddNR91SNjSGIa6W5OIhcp9Kebe/Pe504wE6jk/Mt1GUn82VhtD7
l0Uif+mgfgRNhmsZR3hQml/IWUNXqYQIEpfjjnsgsjy2qT2wMlYwmuchMQYiIKwFTX6JNR73VrUQ
Q6ZjvrEoxNLh+7+ZAQuiAoWE8tbpTvGoSUwMd002tRIKQHrYTGafhRbgZX4X2/iN+GOHrEPSHGqP
6mGmWaKA0aVV3NxX0EtDZhmeSrsvqg2CfXttzI07JkEXvcKkXRh7yynspN3XalW8Le15Pel7p2S0
rbqnGN421QC3O1kdTEx3WuMn9FhHPMw6Ws0dN0G4PID45K02w5AMK6TMWgH/HoSJ26kjf9djdEtR
lVQ/bfr4mlPqDTIHoJjMtlWHIlER5WsnaAkyrSaBBKth4ZctwDApJBmqCVfPdy8N5uX/LeRPxwnY
uS9Cq0jrQv/qUW6U4xXvRjFFzffFPyLfip3IgAzVHcib4ID9jJEEBQ7Csfl6zzljSI8+8lb8QTk3
LMT+UKSbXnFLYxXqaP6IxG1AFCHpsxCxrHQfnm1HFnMyVeUx3de/jF14/HOKJ+FT7pCLbjgQkYMv
WwbgJBiOFpFOyX6dye6e9bvbte+sz5PKw1BlYozoIaCAao0UPdz9so1cmRK/vBucBQS3kCaNN/8w
i9i5WjFmyjWmaKkEQPN3DAmkm8rz/M2ETVVXfMUSXds97XW2c+sRW0A+95j2+j6JBnS43BsVfbUf
OEhkUj5kB3cRcGIpz2T12HPzMo2FwOkFiVRfRuPxxSSewr9GCU6vZWWMWUhPfY4H7FPbwrqlyxTY
vW4i+IgkhAah8A2XtGrpXPPhRVtdE8YF6IrDz44m1soxw3lqwLM5hg8/yr1t4OgfMyjmFI40UiSw
MnuosegMQ7ZynoidF0dtX6NHrDHOox8lWuRmMVeJIfzu3E8oAvXsHUddctI9AbofLu40xI1AjmFF
yYWnUYIt0Khczf+ejizhBJSNMcNX0dLEChksmdF5NUoMgoBYZXK09s0NffWwqb1xOtXy10WCS7fm
bejk44DTeYZEiivN5yg9JOJ7TXSSZXskYDS+JoVDdUEacCAY02ttjjlRaOXUA2+j8r0vUyOACtTd
GBDmFbOqNOR6JH+yw89ttn/soY3LAWbvLVuApddae6w7O+K3k9oPL+KzWI7HCqpQHPi53sZ4QL6j
78rKzRMY9hSmgGCzOJ3bfNA8of2rLANi2N7gZQqIxUI+NLuWatXlQ9ma5npPDIRaatRIqG9czJOQ
9lhazJKlddJCI8AZaml2NLjWc/ZdTsiYrYnad2lgf3wMgyNR4ngnyWqxsGEQBw9LSWTvHa9MX62B
4rHMIXsw59uzPhAMYwtyykDQ7S9nmRaiQ0bp7w0PxdGrcxqyZ5Qi9fgn1j73wAsCBjAxDIb/NVgq
xx3A2Wiy6cnwALbSTOmiKNU61NpPmn0+1QNLrzGyvzxUnHLjpkz7/6CpNUb7ZDdvqgp2u1MGpkRN
QBrYxZziPd+Y/94s3RVdjsDZJRqFub2NzkC39ON8iNe9LWIJjhaNUPlpIxz22ERUz5mbz9ma5qIz
1jOxy30T6C6gL0B8DnPT/XwNZvqIm+vFCsMAIL0P28OR5xTSuro5R6rgRwc00IeVn3eefMrjVU0B
b2D/UVWlwtm1nLI6PxHiRxud40I85ogzJUjHqyiWvz+yCM0vFCgqzqN252XOXp+ymKaubWQzc9nX
MY95RVEMECcodvwLaLRsDxmmqK++E6vsWLr6Zh8xuF2cPCd4Gp7q0BH6B46UwL3NFygmMKSTFVER
WDA4X+L5M7xCF+xp7lBDFjLCxCRq3zcjNaj1lqp90Ywr2vvuaOlfEis/26ASaM30hZqdXl+6QIzq
jL6YuujJIE1FjwhqUcR9vu/iBzJvg+2MtngHiHQmlcdJK5ncLyu9/uKIPMTySaeQ5FymuxIPlSoD
D46L02rVLgu1HYOfkJUe+RrI9gbJk3VgWzUXwgp2V56K04oD2hW4+G8OTBxq4qM/4uzoA25LEFNx
A9omaSKCZ4A9DfHSckokakh4o06vn8Ei6RXVXVP4/0ouuAuZYXAVE9mjm21pXcQBFk7nND3yYfqv
wFRDlfQM0Kk7TnMeKq19saMxEzBT0NbaJ0DySNgQzOTHXGC3SEtuBlZnRCykIV51ekhJ50SfhGMG
cFuJk1J0b3ozkW2ajzqP8mF4D9bkEpu+gTb1wBd1c0RUBmi3WfxyWpJ14PdTWjifffs2q9RXEVvy
MIGerBL1U1bJHvjFrkFLgYMaaDYDYvax7D/BiGpqH6mqLwoNvN/aqxId/GgWVkkCnfuqTb91SHdY
oDh5/3Qzq4XeeDa13AX6mndULKDOt7h9jLHM5mTpoitfUE5iubrtFpFxVbYqwd4ozpUhF/fn1SGV
Soa8uMtdhrWBUIYksZyNJ2dY6hoUAGXv3cO/0c22bf9kyEAzdw02l5s6O8+UaBl466Rmd22MO49n
D6gdqtbOscmVk7zvnDER6lFs6SOlqLwJgNqnfGZyO9R6SBqA+Foi1DPElReL6vUnmn0Dyi3bgzBm
mJt11JlkLSNwgd/wtXEYXGSYFmQ9DXtXWj7gvKP4nu5C7RaS2OhbdlKZXwDexd5kPB04gy74pmzm
3o7oQMGn3/iN25r249GmQSXEq9H/PPGP5Mcbra7LzAXZjAzvZbZbamokrK7g77khx3u9dOVYrX/H
Qz+bh9tyt4ocp1OFCFj7xyxLhPO8uyWO+9dKfHO9jICjwwFF/8z/T7QEg9H5T7hAXjNYYve0XX7f
y7eRDjOCo2e6NAzONWt2hvVuV0l3/WZWVKvWe3krI0gsWxGMwE7kC7yjdMzsK/Z/YAZK47/OqRrA
2f6RYcvOJ3I12f6tUxC/CcmpzlEmIndKJxK5PuUSc9IkfR+uSe7G//UMH+nrWxE/jy5hQW5ayXiM
pUPpCdEYB6mw13o9MK8aBjDpvXhGDWN3SJ3p1a0xegT/t3P29LTMgd4bWgCBltq39Y4h7bJgTnIb
FFSzSG3F7dmRtpIjoB5jvMz3ff97AXwHdwJCpY+8KPxDnkVQKDp5n4mcgQhHqd68Askq+2PKt1qn
Kev/cDla7za1cjbKjq8gVJ9Ss+IhSrG4tHXU2Zev23Kx6+nUyeIaxXUG+nmorgjeJ/fpf5JDd6Ej
C2EPqgh8RWtH3FzeECm1nHg+GabrDJpNC6sItTmjdkCWyf0gzZB08sjaT2bx0Xhr8Qnl168bPula
odoYwzn0B5V3v52m0IdZoHc5v0Bgkb8VjANjoHAXcbh9by1kcHewM5YyKBuy8gK+3ljLyFIDeEx8
fk05NbzIQQhOQ7CBMiqZzMmuA3T+36RNmMa37T1vfr4hA+K5CPJ8BUNPXN1Wsk53AU21kIipXTvy
n5+4oxHWeiiIOF4FrPPyqYnVqz+2jWMHIKQl1wJXSNIraTe3VsgS8B9hhEN9Wd1MJFY5wRX+6yUa
C95k+ujNmJv4KipTkaeO5q97NdyzpvbnLNvROdVdPrwZsO1J/vmc1Vkw0s5HfQBxjU79+DTkBLz6
bg653XdA1qnMbF2AS0YfBgeBhW1/vBXbRRSbVgWlbwkWJ/iEZ3LxlEkk4ja4PY0ZflQ3JQj8Q7FF
cyaXnIlfUUU/x57wDEUafktC91n+UloNHsVHwpOKzlM4oXZvL/TcePMhwEyE66SRs1GAF/RvYYVD
sePiByhcAnOEcKlofZlYslyWfni5MnbyS1gx3iIvWGpuwsbt4i/dy3aKp+5qxdvQhJXZYKMws0PJ
f8vR3FvRSvIsqnLK8osjOrXRyF/h3Hhz5C69gcgoLXZpfiYLeArghRdndTKyPRhb5TQMTAVoo0wR
I62lpLIRV7Ilfc+8DcLMST6JJCGSH7T/S2J1a5K98o1Y2hRSZfpxrxfd17TKAhcUVIYxMkiqlFUN
UCUapEjB58nA3VD8z+mWAQVf/AW7EIXpCY4nnXSKt5zVctKrOhs3RFU5RHaHVMKfMt1uZ6SG3oyc
2FaBnd5Nde2qchwbnbBZuztvH5eUxiRuhGS6ZDwplBnebmaUMlKoKYRldhhOvBf5c4ja5v/tgKab
sJKQdBksg+aQ5Kormso/WTFCI26+SiA5aRHG4L662S6qk8GgEDw5IxCnQ1kX2flHqnrseNxFEj2w
nNKljpvS6upSpdfcBPg0YDdNZuzWjN3MCBmhlJY4S1f4euYH+wiI74X5UeAwDOrcBQWLeEUWI52Y
38JCOgce1RFWXFNXES2P+n6VdFmbQsx8Dv3zQj1w5Ktj9tnfZDjwCFb0bPgGN6CFq0oOYgy9m/S3
AopVzIPjP3OLRJpvJMRFnA4+2NaOjFVCFkC+7Ds8cstR65fiyzZVtqhM2yJSkZggM1Ge2yI9obET
PBtM0h++NufJZLJdmD7piMduLhKlSaX2ODYvQPeInsux7AEtM4mhtA1d2O7VVTL93XHp71xK0W6s
1nAlL4dN93f+gjyV9s4ZmYHVxu5WFtr4k4cepGXUiVQB+I64yKWihzUXOk0qClBhiLF+rB3bPYDO
OcfiX5nxLicZm6oeKrSkaImURa1WCAVe9q4adP99omFPcBNunRKwzeGAHnCcrvqz9699FcLupJfb
vdhBT8jOyHEZ0LuDlS2Lc/3R6LtpPhYSl40X/Amds5YDPcSr2Fhge5zenOm3jz94a/X92cqDcYpe
mdRV3C/DQKUPD4JgSKfTArrnPHN4x+4Y5ziuvljEPdt7DFmUfGsSiIcpMt04FOFCYxo+w+Xidg0Q
dvoe0DYmW8OQC2Ib5Wmss919gQCjhnOwXbZqdd3mMmHwDEjr3muOWhcP6XoubNbmDCMHdLvYQ7MY
AkvZFwCTdQom/d0tbUju9Fvh54Letjjcie+WRm9YNfM7IMnPepgjFGbymjW0x7QyKbCLxd8bypWM
zDw4Vo3U1DLzejVf7XVIJtoS7LSDxPJf2G5V9/BExnW/C8enWVmFk0Nr+mmkO+iEeNV07CyBmkNL
cH2rev489gDYxuaGBwGWY5JE1KnHXxTSy8IQ+6iWUXw7XB6qd0/u535jB7Hm4dTn1UmSZqUTpbO0
qqO0Z3tCjdlwejZQAi5+u89bLSa2qM0ZWSJG7hqayzJfJFCBWJI4YRw3Y+oaxSjGkp2hm5SAizYx
7vB9wc9pxPU2gWYHxA9e1QK0u+OVtrXAoCAUhf7jcLy5NKHdfUgB2r9j19YJ3KCDGUdUfaJb8k5C
S945GChMp4lkOHf8zTz3pXB3EQTycwSojxju14vgQraQ/kK79I7UOWFRVwZeZwnd9ooV1UDAHQrw
f+KLrWUXANsT4i1onVOBbPVtDVnaZCpvxqhXTNJtNOkBVvPdCI/8wirX86Yz30mZy1GHYWmBHVSJ
dTsCM6h7mUxypzzwuJKDTXry2vyI6tumuNn1y5EThImUHdASZmrZWPHX3l6OUyz2Qs3WzOKc4678
YQ0JxajfM+4qb2+oPOcaEnav5P/Vkk5rK1DZsiMn/REZiI97Acy6tDtPl+A2ArRu9oS799wxtidi
5QKhrvPLRGF7oqdoJwb7k1XlqXhDXLH0zk1NBBPRvogaGrpfTpMPO9eL/NTII4I7truEM7BbFDgz
fvq6cZFCOkHVHMO0OhTI9yjqAbTc9KenJR/K4yKv8z2c7U3SHe9OcG/khOH/1L1aaOBp4qfs6G+0
tiG5HawDeLRe9PKrtX/MGxCoh7al3v3wPczsTyY7aYzakjOxFp13ac4RonZy3EJsaSzLreBqYg8e
wa+X4HRNrPK7e/AMBMO4VE0DinXjEloTAfnE6zyahvg9i8ROjMVdNEg8ERO7JYZFVVamiPwEKV9+
fQ2Y9axj5XOgi+LOtacpB53Mp9WqNyb/tLZGVVHt869EtwtBa6X/ykrFo1uzR202ydIa5tvp+VUN
yJrwlvYMQCoSqoyd4C7EZOL3yo42yG+fukpRpI3Ky2m4NKcJgWWHX7tC/Y4E0Zo5mZ+eDKXQ3UyL
PZy1rsPZtAoFRKhQWSY0XDTJ4/mP8Mvi05lQnEyTcX0rP5OOFoKRFoSHM+Ow+SPkXQI4a9gZjlYx
O/Kj72haA97nD1ghvxU+1nCGRIVDQOecyu8bjAQy6i9V9b/2yeekCrpC/NcQjm9u32tSNE2kDPZG
CMWvdCMO6d+VNFeS98qc6T0hI6OiJ04ttK+hA80hUBp9GUeuaCbR1n2KVYcSYCgJo1Tb4hF1wEqH
+GhcS2lmXPcsYvGdFa/gSGr2qYiEGmWPp/b/Ln9X+OXbWhakpS3n8xCKDtiSed3l2q39s/9ABdAf
+VikYK/f881L98TaqxU3Jakr1qO5Etaq3LWCstXy0wXxN4BLgt5xhCOPKWU4kDrVoHvT7Fjri9CW
LWVANn3Lfr48bmnHjKIuWKq1XaFF3PHbyzPUnxG6L1RjsXCi8mUoVUoPqp6HrVZTY3WqkRGIamWd
xqOseB5Z5mYhIalTN1w+iaGm1cVpjaPpRIBMjniDjB7EOhiXcC5q2FK0GAAmpgi5/A+gLKF0d1xz
W+OnEUpmCNp17ZdOohKYrY082nvJZOvlekBqZkhMZ0ZjxI1u/eRg5CSskmgMowI0tqgJXlsCVnmY
14AC1O+9bTXnMkEE+6NayaaFI+CXofw3OlXvAmooMqyURyXOnU+tO6HlhHuDgMoLIoRh5u/nus3q
hUOjzkCcbeaB/5b059LYKKlLXdsCr9aTwga4Nx13uUKaNx/duU06DA/BUo92Wr8mmLn2wgLVGiXU
9E9UBQ44vFjB7DqD0zBjiDh+dueMpMz5MkQcbZzAB79mEbZ6Syptfu1JTsDP8LluDc/EgdA4C1MW
L6s+MTMmtblnplbzScZGf2x2D1yd/LyW1uAzHym3AL3aU0ESXxsGHrVTKnZzHqqVMWTl8jx/+VT6
WubrrAhAIU7repMMFpbi4KMSGgBx+0xKhGCOOhJD9SqUGQ/TlhJ5pGcegosLu+BC+jXoiNWUJxnn
pwzMduZS06WpkwvsqWTCkozRQMUd4JxggZ2TKoH+56g2aKEi5Mz3FVITXNhJh3umhFgcN5/rxarB
YAnuh887gD2d80LbwDbDT9JX0XEiyEK7sF+TWgHa5lMUaKrz2AfHIScPNg9fWTRrCzVek3aCSTM4
MB7SwtHRIkG0zCkVL1sEhrch0b0LKHWKU14QNCmi2yCTCCzYOdmVFHjPraQQShYk5i44kW08llgP
2TBj3x0HrqwYkXRFnwhW/obriLdyDx5jUXf8GzdYAdpbtivIzTSYHOQ098ziTiLim7zYk6+MyGBS
bBsNgh3GKmMwnAX9GX425kJOFn1T/qg+zoBWrDEULHgDebPo6vkm5++wTNutcH/tzYMt2Yer52PX
BA3Zg4JswV62hHLah+G1o2pcUpi1PfSvbjj7To2y4mlfNV2jryW7m01mZJasHDISJOs2Qy8ROKpC
MNe30Kl9Eo/ME3s/H5n5OZ+RSR7KHugqDxFWhIFta24Y8hTZrXgkCmQa9PVFmkjzcn5R9sJvQOrH
nHFlDeVEJIXhUmyCIq8B84wG8aJC+0vsLpBl6Qe8DWSDEaLgiyKf6GsXUYOh8ky7nSTTWHcRpJ0M
22cIrQR34G7/jZ3emQTSeHtw4CyoH/3fgiIURucD/28UUlL79vSxXE/ixxUdU2Om/WmiBqexigD4
qAtxKs4jL/tDPmusYrhRnwKRlpQlb7BlybLR2ho1PALaew7eFf8q1o3t/iTKC95V7Ja+//WKZ9CC
UJVId6wY0Vjjmj2TF+GHdul3EYlAptpP5wy/IZwU2iVhgirJdJag8M+/glhHjzYWc2M2a1nBH84W
j4tM68hLVvhIleZCeFxZS5r9b9ciADo07ry5wyM63rtSI7IL/El34mw+z1aE2wfvsvT8CpuzcLBv
FRHyg0qyUcLaxSVwaJPNCnRUyZf9XrEcfEMMPZUZZ1PBdg0fOphq5qF5EhqHvfrwzABDH/B1FOWV
cRKZgTVTEIa9jZ5JqradKAabrFttQ51ZQojXsu9NXXK+zlCQJqAwbxo03IMDpsg6MOW5e19iFHw6
IMehe2yXTxSeUhnemc2eSuy9wnfIUtTOi7P8L4ziuvOoUTX0rtUGswBO3J5wO47cFJCTXwFohGGi
H145BLKB3cVYGGvPgVNhufluNZFXFQW3WG3iG/xasJPJGAwY0gGHC1FuSUkqNr1/JJqnzAXJzu5J
DRS9gjOxFNXpanK3rq7CeTaNrLbUMy6uAs8QklwhtmJtPG+ySGvJFxXlC+Lt/S6Py5bZ3OmLWvy0
CF3iyN/wSJdhE6/TXE5sAlnQOalbgj8zFuMiyQX5KhgzVu/SsOCtY+mRoMy7QQP1PPcCjYhNYrHE
VsM05x9Zb7zuUSDQSLlMJIXFicZsOLV4lFZIiq6pPkV37fzKbCYLE9/7nqcAC1Fljwnf/e8Nn1V2
bTvZB6GoYt5Q3iRcxzAi8RbvaGgUR7x+DqJmfsinewLKFnmfC4WZ3uxfag+fktps+eTN2QAqPdB8
7owBgnKnR7he/2Ds4F3NqQb9fLvP3je/XrxXuuwsklsWXvnk31nnEtYVDAADmpOVuI3FgzlFTIvk
nFn/EXFJgPgT8V6Opu04gX46DZfPs8OAq8Dd/QyypM9IE0chxxoktC3WaWrcowVUlNVqgLR+4MhG
kEMW1YfYc/fuRIfnfXraL77LWjoMc0MtqeMbdv8U19YNS0OCnQzVfDjA7B8KIQOh1njBx82ofMlh
DNwcdAC3uK7I5MSCnmAnGJ3CnpQkDmWgHH6KC+z0ImO3mzWiYi+ouTeg1cHym0UkZltv2+dIUakj
QqNdURyyaSej6NbxhcbjGw8vy4y9OWOso1jCk+S1PHBcMqyubWMHkppbhjdHY0YHZjZBu9b+Nn7z
xF0vG8w2cqKH9FRqBs8awFlmgARg9pgfh6nWYLEikghPlht3vDW59jwax/n+2I7rw0gv4dCmS9bF
30ehmxzn++4QtSZTB7hQ2R5wBdXLPg3ZLJNkAj+kyZsAb+xeDlXjRbKJsgyXga1j8Y+g3N/EDyhB
OiBsHQ1Oy4Bgki23YdV2gIxovArOF9owIQGbNhJUovKI+OnIwNjCJmQHRWRAcPXZHoj+otVVyDp/
UyYRIGTgYJdXdTminGVHDufqePeg2HSYoTWV7Ujgratb7EpgRfQz/pzaZiYVU3RI9Ntewk7wEkOB
XBTmotBMAGPnyd5hsacpxhvjN4kWxkqJV1CGFCG3nqe93dtqbudBOas+ClFdOJZM4sfOZ+ROf8mt
0oCbmfK6IZLy/J2xyZ0CXjd87pwWQ/EEI9yJfxlovqMYqyOyHOFCb9VfI9vvcGC/7J+S+i+d8HD6
kfr17q4JyDxhBBShEznEry6sQVfOrmrGeaYm1AWyGEZ7p1oLGcU/B5GmIUVRj38A0oi+1dwiNppH
07ne7RPO1PqcuXw+8MEg7BjEZ168wMEHdX65+NL/YN30oUXAcHM99467eaHPsBZ/8TZUbbEBUvPU
rKt9479yshX3LyeRLM83txbLlPTImEUh6d/4q2650advuitN+9HgMTpFryhA5dw+9R8Vp/tVubWS
WVNFOqHBNHUH/qoTMNHaKbx+/DHOLMOvqbVm8MU17Jkdik35TIyLx1+kcHxyIVjxmE1dNj/Zp5PV
ZvRfTLJJ8dg4wyV5utA8HOZzEUoDo/Kr52iCAOSbpuk0fq5QRUaN9LiUyGYTEH4uvAKCfgLVRmoL
GPhoY3ytq1CzLuAEk2xs4ZC7yYO0xZipZSQYbkk3No37VWIZEAi6F6LBSTMjKF0yZdfWwiFeggUW
83TdPiRLuTQmm3yFnzlxtBPKrj/IQjtfMXrYhZA2taV4fW+S81BewKmsVwK72c7Kfym5KrFuX7yW
N56mUPzP4nqtbclj2r7PE+/BKwL8N8H8j+T83aaSSo1RMeXB5n8BzxqAYuSCV002eV1zxHon/fd3
JtQoUo9M1KxaAKJQT0QGCOMllXvxIWG3PEa8NDh4IKbkRUAeVZNBjJFDnSEWiIpCQCehx09RHG3O
NQrZP6/nIn5KRrCvkDrFJrzHYT7NEQPwBHCzKxwJKAgeZfgDSkDKvnI/1W/Z1mz7ki+ekZImXQ9z
4tDlYssdSoUA5tntktgEI9X9xaUkj17Y6ecYcfl7CKjdd0mAXlq1OZJm3XlrbZ25cxybpqoRtm6F
lbnrXj8SlSBZzPDt/sT6Bi1yZtvEJE+aM9+ejycx9nNAiZYzqPg5vHlJdrOpzVLnLaQFP6xsvyil
0ndIv2oYWwTYQ8jcAKIrWk/CdnXp/R7ACnA4gozBS19JRGMKbWf73oxJtESVBStIu50wwBIoG/Bn
co7tgryCLWTXxDUp6Vkdms09g/1Tje1psMEd5ufykEW7/i7IuIj6E5Fvs8CLAdN2Z6W1kMBJ0zD2
9xC5DGe1ujZqtfwDIKCLp8v342+zHivxaYfRSnFsUyDD9ZK1etyEvM5d7zAr+FxOtNjK+o4hv0wC
cdIVBxI2IeHQzNeSrD5rEginlseGgQS+vKmt6UMyZjfG00o3RT4HWpcDSj7l2WIbQx0HOTzbT9SQ
ln0K4kaBREpSB3/jYhlqPLbuaYOSwjwk3NqpcFeqBhEuJgJYSpuEeMgZM7OHcquZGHWGh3/kZS6U
kZh3G4jIMVywXZtCnDhg+EMazlFPN7uPm47N5yNxDAXx5Uk6hAozjyZqAbmDIL857CrNEINWUKk3
1IDEtofVsLNJkKGeiFOvNiA1ysHufn1XStEVrjlmZnBAYkgJrZHVVUFqKwel46i6MY15jMP57y1j
2qm3QysMOL55z0EXbi22qdYWoGQ8HA0mECntAeKrIaFRnaTexOXy9J5YlARQgw6YcSw3AafdoHa/
Y+zPMW8FdYkaWjoUBbuEAwbW6CZwSATlRNAMNzxvx5ToEKEGjx4Cw4ei96hClyrFHW93IZgyH1B2
3ntU3W3Lhu2a9fGU5+i4esunDXQUamzjQVncxqArttarkKAtWVQOSpMEAf6Uyjs5zUJBcFZ0w1zr
GW6e1Z9kZN+AKrT1S+ujCvZrutvUsEs4x74glJ+rMDt1Ht2JBX6j5NlvMeC0tJC+GZvEQj9ueHt7
l+qzcWeXTLC4syHT9fiumX891bdQ4o0KL6L8GPVPbp7JcLCq/pnheDT4jrh9vVjPk7Rv4oA6t20S
ykrLRj6PRU44F2jp5g+JFCNx+1at2O4dkP+/N7PAJvTposLJ1xXKubZAvx8dC+S7MAwuoMBIXMah
7n9V38t3jrM9AUporrtZrkGXI6160HPQEm/L7/9Jm9VXh3tF00ylQ3TY/Xk5gWTi7aC5bRbizEsE
HcSMRJawdkJ1EZVdlp/KbmX5/2NIpioKd6x7YgKLBu9lwybjE4c+CvLGkD8jY4wOBRy/UjRwa554
/WAWvCWvgkvsDXBwvL5g+t1/TaJxzg7+0ls8ov7DTd33ISHtseni9XIm+ufpSh/y9b/nlAxWUOPY
pM7Z3C3vvJIdkpBtXPm3fLFzNw9DA0rb1ZUpcZgASnIUbYFQ6qpktGNHEzHeCeVKLucyRNh+wYCo
FaTQEZ6sjpglZ13eKizC33Cjz+gYDtEh7uCZYeV7vpl/BAMzffi+WrR0roroSkR6tobOkvuW3jdn
MyC1FlzjxZ66301qAMJfrChFGn8eEouthTE2+DZWrm9/sHQ30GXMzzWKCe6MFs6YnlatVEu7NoDP
7uF1FJd/BfFicHyKj26+iuDP9p3WduFL757Jwjcg32nqZwukfUEfnriF82giyMV1PCBJkqPL/t//
H3pXIBOxF9OJUfoA7uYdkJx4U4TxY6k6G1/ltLzJ8jsejyWyno2qC7Gc3gPEbZwDS/tcBfPyT69I
g3dQlhxl1i8a3FnNxKEJbbr2LaXHNexyoaI5sGfme3bZ1UtXNE8M2L8UMtpfKsrsEct1YoObQnCp
GG73yR+8blzZI7XTmTo5vogpigqb9XYkIUT9B2iaQtMbM3q8FLoNgRadRQ/81v9UsK4XlhEhsj7D
A4yGmKaPYTSb+asAg5JM2P+0H1wyhtgBRUrPeYGOUjxPmNW1hpZwBvlH2Jm6q2nMieI9cNcn3aiP
X7bQcZCvLSgvIKCQ14uIaolhPCp8cZiGQAV9gF8D+qWV5HVf9A5rZ1jUI/kKHovQswBkjfcGHExd
SUiX0L+W5T+JbRrIQQdcQGryO/S5lSIEedz4xosXXttBvX81eQoXcUjzDRqgR2GNJ0gmhI8Xk+6S
4tLYKFWetCY/CMNJnd5VnC7XmJzoNFM6KcYmHFWnmmDHDcpOSlSIqy2vKj84vrj4NxXyqStPNGSU
FX9ohFnlA53luUb/3UejppbNm/hNgLBjyQ0mpBIwmD658sNkglKlv5XNikLg6R/oNSVBQcceORAk
n7DR0VQUQ0horattiGaK9er0if9fI1eiZkD5xqdvy3BjHlCZhAvBxcse4IZV2/agUzn/PSI+OGsJ
QlpCzzKtkoJLytnXVjhNL7OgM1+kYshS/qCJqZRbT8uRyA7YXfHiQS2UF8XKWnGgv7x7y/2aYkSX
8b6omPJj4gibLQds/KG4N5Vsr42Eq32FdHIfcng8CMljg2JOEhWMAKnDIAUB9tSiRTE2nZjfS+/1
yHJwc2Hp6QB6ySA95aCtFSZCeTspgnqbv4eOCqYnxY6ZCWGQD44SZz4ds6pzMy3DUtynt/3z9qwk
zRyQdTrnEo1+jjdaITzEMqrL+2PM/osB1UGVrgvnbGIg1zaHPuU98mzy3bZ9xS8omoVCr9FuNwxF
PmQk1VC5pU5boewY7thk5RZ6+ozD9OOu11RU0+uRlOdhT3rwLQDUN2NgdjqEfvACG4uk0AzD3dAW
3WcDBjZIta7Zth0ZQdJ+Clb40e2I2myt9ZgultlmtYYCSqF8OKORf1r3uPp33rcellrPH4fTJIrY
A5bpembr3QMc1o5XwQRwgrBt37ZbEIuSbM1NwT0zm+u3tm4tsDWs6+uMGF0vQtxckILGXKb603jK
CPSUm9OqRhqQR6d36OmQc9cwhhyCnoIZHrbSMQ68dXIISccE3hkNHt5sL5L5s+r2a/DDMhihfeQd
oa5mhNRhbIwOMxFnsELK/Pr+siJxuQmgpOzGdwGR464ocncQyZOU/ggYpvuI/mpshBUE0bUoX1cl
3jzJEAK5SP1/7PueopsqwzSodZd2YNc0jKY/3q/lrc3KOO0yqiRFDehYVasrlXjCFJmfsPTCgri4
YYgal/B4tbxs1KG/2PentXdrlIGxFA88soKesAYW+9uwxXboIPdT+xEgQ+BRr3j3qbxqX5+f1Sz4
5l0na1JG46VduySqNyjMZNZP/IlqhUcN9vMbahNYj2tEI7wfPvXgAI9gL3lsRVcThN7MNTF8u95+
sJNGt6SBQpHFzvsMFgN0dElKN37eCpS6dA94275KNwfyMRIQt6ryOZ1lEOOarJuZCDDWxKCwsJvd
pJlLtCrlbOFr4DR6uztSP3KAkErt4XEkCJnmTAN58qpquPWH7OOmHguNK6vGGnwxMtmLmQKIqghz
78K1Bg2musRB+JDAEgKxt5npS5oud1t/xHrDB64xQRrUISBOwOD6J30WpqsKFmdmyknvXpmxY80s
3wHpexJMxhNA9ja+2iPzSpPSaos/fd9YGf4mqybV2xI3kKA7+ZbDRb//CycaCM1ZObhUEYdqhxb9
YV+TFhOqjHGT7gzzB/tJX+mJ5Rn7IvlL2aszE9dgdO3hWoLcKIvcLUg6VOqCLqxQ/UK4+hoZckHl
fOkhdOHJw1D4GNhaJ3aZh2vm5zVh7UHl2q0zDz6P9jX7ekxyMs6NYiVZjJWxzK0G6uxGus3Zl5Cq
0tp2bTRAMqpprdIzJ+G4OEdit7iotnaom7GVyNKzd3K/UmZhyLxwgpSAKX6yLuIrZIAltES+SSvK
YG9m3nAIfsTSaN9UsDb/TL5WVpWMRx0m+c9t9x3PfTNBQ7KlPl8DNIM5FAeYVKlVsQUomCtZtE5n
OfjqJxaSAn5HqlX12mGN3/2BZbWJaSD3hTstQKSUQGvRpJP7WjyAFS/7F+f2lzTdYAC44tdYB646
/T5zUWbekd9LvMNDCypiPw1I4jOuQ4Y3d/Pk1TpLaOyZV7TDilnw/YUS3bpWXrQj3nKJPQeKKRXs
UEczp8B2tpw14nk6g8JVO8IqMGwGJJhFvJuVM0iWliE+/Uu0thTvcgln5Qs3l9xHLfpH0Hglshc4
M6Vl++DhcmVujNGnxUFvs7b/QlJ8iZt8AkNP88dsvcw4tqgsA6SYZZIhvEPXOe/E6qE/RUASoIUq
IXN1fDK0GgdaTPzTFx6BxW5qZr0eQ53XvN0WS+Y8HR9BZy9NnHjbTzUwiKAQSs5xgJI+fyuQ6sSa
5MfJN22bbUtedFUAsV2drjw4O53/b4JEGwyTakwI0VJSGr1dd1t6rQ+cE6YNCgyPCxx9EotQx/fu
OqCgj40WfXGyPiupiboc8/rvluAKbGYYB9RsvfS4LVcCt0Y8F5thoEV1vzNZ4vH3MEeZrqGY8Cqx
5fLZHRG/MWOdSHe5WBYCxeoEF+qRBxm8S/1QD1LQZNjbUb4V8gYpQbER/rkqwNQinE8vlmeSSQdW
4hXFmCKug02SednIVzVhW4OFrXdD+CaDjRLs7VoXPJIbTZYAyd7pe9gqn8XXOOSmF0xNrmzpYxFp
o6uFTZqz6up+V+j3Bke7PJ3Ud8d3eAsmkjbhWqHZczuqpJixoTCVNRKPA2WVmbqGlJ3yOUkf5v3H
RGJf9c7xOY0QzFgRfpNQ/SrPn7t0HT5QnbUxeo2fQ3eKbcqj1UUhlJ9WmeODncIjdsArPOiL14OR
aSHf7xYWBLZ0O6f5bgIxHAsLcqpFbb3Bm7X031DkLUPJfkMFRukaIQLTbdM0xpnhNEuf+UiOpNwk
gz4gkoBbW10AuwJyBf3u9Sc8skAmzHlHro3aHM/fFCVsG0j0PBgrgJrHOJdvfpQNuWDL5vME/Sju
lh5XIgUGqQBF5xNUAH1t0HTcXvlZE3vx81F9hN5VohhwiB2oVDRApYmn8oEk7jsIO6nH5qN48SNU
QthaGh5jVdi+wwx3+VW92EoTaiqeR3vO99iXSsQ8hPedeehG+KvIsFowpFJHrWP2MoazAhx8ZmFN
9jMtJ4TdtyqZ1D8kjBa/tR0DmgOFH2mk7UtvP4ME9V7StNnSLoQ3ZH96DkuW+KZjrQMNohXXOaOx
xXb05kCT88Kb2I5NFCVgbpn+3Ovi72jskev+6UhcnBTfGfb7MuTpQpi9D+REqrMTszqlPDfgfsVJ
2mTTOVCSLL/uLIxAfQzIIP6Xfymz1osn8w78GRWEa4o3J/jt/oCyBgcrbk/c+ioL8JqytSCffHT0
vT9lKtnu4lF/M77XDhVAOwG+Qwqqe93wOFR3CYxtB1PE9Lko6RPSl/Gf14GYUXenNLyZ1aUp+Ndi
BUAF5huY8RkZL3SyGYZi7iHtsKzQ3bCkPHceDmzwxvTGhwxf0/+NfkZ4St2ORSCL+740CAHIbVhC
bsxxqY5/Wi9Oa/JLfXOoo5X7TRIEEzFSBXs7lnBzLPtAgu3oeuJk0iqTslM7PdYdRrtvMa5pVhIG
SE0OIbUQ4RDxlKp3x3Wmk13MR1h+ElZ05hoq9DFx2tz7WVgckD+6s1Ul73izNWbusMhIESg5Lt6q
c60oyaH3YtT050oHM0ErvZCwm9VwukG0M2xavcBH6U7I+kvPdodzBW6AC3loyFg8oMDNogSgsJee
7OzGjsDjxtxEs/YKTzQLGCfgoNcDNtPgEVeBpVwSOYBwgkvYdGaD2MmHtBybykkQGQCFMH0x1g2q
CR6XXARy3SDy9+j1TS2BQ6re8ztFh1BzZexiWdGayUdjXqY+BSg6drXziJpZq9km9QrPx8WvtNfH
Cp28UeDG+gv/BLaBApUNs15oaVr5r/pXX17yjPtg5o8ri1y7lV2vpGakjSMaRojiCzEtjPqwE4fa
T8ELPKhE4TZ41XCxBFamFaDXZ4s9VPCdyKFaoK9GxeqnMaJFRzzzogo6g/E4L9QX4iSeeVRvQ9hM
OMg71Np61cwzwsgXFGeiQFKa/KU+IVh3kVEmN0fs5vclksfLTKc57BkjDoJtfZwcs9SzEj17Zpem
zCY4L2CMF1D9rSQGiTDbShPeEfHmxVX1MsXnxfYQqsccWG6CP1sQTTr+XdwzlzLxvxYnlUAZd9QS
P1Qr4PHU3xuTStUVvFkuaAt3InlRsTXPa3+Qu8yQ5kiHve+g+TLxzcpo86j/4VGlxZ0lVPLwce9x
vlEtGcQpHwWU97irgnt/pYrzgA/u8em6qKX5WTCHMlXGpbK3zUyyvtAloPYfJqlDQUMEHMsInF1Y
xSqO6raAyquFTKt5pBEvoxNh7nKLorJE6a4APC/6DMSdBwLfJgtUMtwLtdpNCcmFICKeChoVrJKR
G38UCW5rvdt0Gdn4Bc2Spz5yU4BxSYTQXnO3ZPieM3FtHa3AjahoGW7sjFCNPAs/IoCmPaQy+jux
gnUuJkm6j85PcPHZDEtzCJOY5XQCUUT3gCqzmWFjOxHetF9vRUjqJk56GDN29pohA/D3TO9ohgZ4
U3X0+fAJT31B05p9bzJPOc2BG7HgZBGfmecIvBoIGNmCjz40fYughQuuCfdspVW5FtyEHAMo2Q6i
AstGZwB7bBG/TsUHlo816CfuDGJ7bJsTzK59yyQEFPAknUj8FTaP+1fHgXA0WOuXDoFDmBaxQFkt
88bWzvu4YEH25bOKBKP/UvOmo/u3XtQAu1eZWx7zw75fs4Fx0fSNU9ZHkQkUicfbkSmRd6cOUUjM
9DWdW/PHJCKia2kR1ycqQ8dYAdm5bUHk6JWa3qyGVsxdPpvpGnOeDnbxEvAqd+IaSqJku/Re5f1g
gQsktI2zMRpoPVy7GcDNBbF2OrqN6p0HCjPl64tBPWRQ2ALXDuhxUiPlRPijdyfe84Eycn39rxfE
SWEKChc9iC8FJLMxMJQRlz0S+ssd+/SFrCH1lzC347c6p29e8XldvqT4GvtChEdn3nm/zneiIXVl
wjs2Qm7TBdjp3tdaU1KeSlapXSqHbQBY9uBvlz7DPBzIp0aCu5WVBaK8dT9BI4l6em0SYcXTUCEk
9j0hMYJAAou4G2unJRdi8gb2J9Nya66YmTQpYLz6P+4CTHQLZh5fxf5qpyXiNNzZF6GGWOl+LlTy
nOIuVSXLTuQDkqyUXWOWGA3JCOGmTy9VF2cqA+/LpGiLZbHext4Oe5i2YcWzykLTuQ4NbHXeEVXZ
CL0o6LOibdvjIJytOPJmYERhRE3hjZ5bsnnY+mKvGe+HqqzujK6f4HvfDcPKu9dzYADfdeo2Jd5a
ce8Nn2v5Gs3p5pjRa5B15NfLv+79WY80hnyl+3NVUN1nVLHHKTQQryLlMglz0TbnlTlHbuGtmBdZ
vzs+KReBO1nEE10iW1nYPiHMI4UzUkpG34WXLrRXCqVPk2l8d8OPW0k5H0Q1Bqi2S9eddYWy3vR+
NP+d/C5Egw7Ciyu3SydMJr1GuiHh29KIThjBZRebU8MY/jq5+Y9fNRCggYykpkcWMc+MsGHaDyx9
h189U0dni085SB4GlNlnpPRUzxE8jJAhsepMMRVTJ3Nhnkw65ptpRvkSmtHFm8NpENyyDEjMHI0S
ezI5p4ukKbFqzeOLlq2ULOROJWvY0wQWSDW4qAhvxAGgMj339yi0gRyRyxIzwQObi5qQfteIH4qV
yOasokPXa8yCZzBGFJVhB2yFoKOuSK3FM7bLmN9BcglxyVWBQ+HfS3MaaxuZaa8n3m8NA7RXJBK7
WbRA6RCq5njWVBiQmONlsVi7QtROeUI8+iw+IYkdkw4sWWwpxw6G+Y042xmAORXxLD/IRkOlvaBl
vniqEXadqIqMT/FtXA1dDS5vNp6365SrrbUJaS+eKUAwZZxKyyIy4N/MDBQcuYCT5JaA57WymCR9
biN4GvPK4DU5sr7tscJ+TycTXld2huLBgOkZsiWL9C5O8LG/4jkG2zsdO5xdr3ZF/gSEAUvjLfHw
IJ/mjLUf/feK4Ki3G46G+rFnpKoK3f3oOITm0VCgOFdN6YWKHhUKigfBcseDLLIDYu+zV7zQBQIH
D5MfxTgz92t2LY5+O2knAtH7xCVpfcgmxeYFxQiYgp9KeDjvGrLfzxSgP5r5a1KI1gkvPmWYh7iD
sWGtkbRm9lPe0jFiXoAKDmrJKUfAsWcsXDZhNJ5GRBp3ZlvIBs45+2t4rXcm9KGB+7beHWUvsdfp
k0qapL7bYunkiwQFPrr3+lagoDPebB9VhhyBHSf2r7qZIb/RPi8iDqzAYkpC3T8XKXOS1V3ZwGVM
b7bWwvU2cPjWiEf4XeVJrroPdwyU4BwcLk0KGIrtmRQRv3ajV18cv+xrzjfB1SWB2vZbuQYGFXc7
0oTMZue2zBM/GmMNc6Zwd0FMu0DZ1Ce4Fr3GFQa3AzT9/vc/8WrNTjyQaEqx5gUphcuqF5ZlWFEh
bEgA7sQRP4MunILYR5TXYed6MRClT2fS2H/Bjf4X0zCKXkhmPEpxY0JLzaziZMvX4PSdFBeo+8MJ
rYc01AplQgHasD+cpTsfAKifyzau4tTk8PIba53wL+OBB3b1CBIC38/uPwivvogtR/oBgKNQRTyh
y6YU0G5cA0lQ55rTfE9OUZsMVWDJVXyZ27xwQh7Ww/vXLZbh1zR9Tdt8xEj2Quv4/iJm8wBWz10t
Scd1m6U3ebcwqM1kGuPHauHRRwwb1XNRE67vcYI+0SflHWYhKI7w0xtDkjlWB9qKVSAre+jEy9oc
pLQ++75oAaJNMWDaNoJ+OE52ryMC1R6y9kf4reoFhFJKqXOvOo/moDrPdHmJ1tfl5ykOfYJZdDkj
NHRM9AI15dceSvQtdL17SN1WPmKfcy/x7bxVEnOjfw1KWRxFnIwbLbAZKLTQqVQoEn1HHveDbSNk
owlMCzBDpqQ7+c0N9xvAJJrXpxPYPoEaXfYEUIcw+AgJs3vVP22S2Gjnpvx9mBZNvvJqOtw0C1FB
WCajnTck7ErbCPTnc4bhg0SQ4rVEMpAw+pe8sowXJ5/ZWktyetDarXLJ3gNS0aarV2mpRsHrOSov
QpQG29o3fZ8XOvnHZsrnr/zwsZlR4PueHny4dwLusKP3PC4MGlXFW+vLI2blWBAE86rZU0M/k3r+
ruHuzDXmQ5rZg6Oj1kK6t0Mh7521WzXR/zxjnlzbcGiWSY4LseYp7+H97bZOFv9Mh7ZVJ6FZg0no
lfQFMy2u+Ldxt53ECCMF6bzpvYes4SdPlCNSdxD4Z2gO+E6fww7D2sRJsollNoIFqGD685aN1g6O
nQelQBLPj19ODLVk6+O3lxIXJrOgJbbxW5HnEAHJHp7EI6ToWji4LUto9OArMV5kPbWxTYGLLBZv
EWHKVAWSnz63xcptl9yiQeAFyM/t3G5YuUjHYGGEvW5eU6M6KJCVU6cxP3ov2ySPAzvw+GFo0gai
b5jIioVmZ+ybFKSwATVPJKiyMpXUCEeLDzYVym/PfeUuAzeROrFKQedknL2OikeziaIcVvBgXFfk
Ua/Us/fbGa26Inzk16jORTLIPo4WH2TXK+CXH9pCznvyiNCWxcx52p2xkcAScZFpczi8dCOZ28cV
BTyn+8nQ9qYBPCB1bawmtgUqcqgQRPMW0CtuxfvDwpMFYMNkwC0a4uxkt5hmNQPpDoBNvfUzGRRk
199jVIDrciSsMpakcpv8jlP89u3Qo0501i5YoR+0tDpNgI2iPxHwyiaIb1MBSsRo/89NhG+s9RIZ
OtNAI8rs1UZ/2XxWucF3phmc5XLE/HjbHrm1cMaQg5w2ZYcVEZEmlQI/FaAxRicGTNf+XeneXsOe
7ezin53QV0pTMY+2dr3IolkbSnUngXLuypb9mtxlEo2GgVixdlvnUgM4j+sIPhZbknN0oAMrcwTx
LJTjvVup13xqUuadfQZOMv93cpasoJ7hUAhlpEgtvWy5reUEc5yETlLkF+yML0UiycpSLz5F1vWN
/7dxhP6Qg23MHAm8HPLvKe/lFbvzBd7xjeotQVgu/2USOmEclZOC88jZ7kRLVKmpgOJestCe9xy6
TjXXuro6WeIckTGdABhjpmeRIH7CsXppwXJWQRdr/CYvZz0d+gH86Hi4fi82tah48boBKp4q0muT
EBzKHckrcnTTg5kBbin0NH5OU+FUsc+Exy3ezBLWm4X99zZdxOMogsvTnkNd2e8f4Z5acjK3wk1H
iAaHP32B5zrMTYeQORPxeikgX10IgVqf0EsLtqtwcj5hI6k0L0KxB1yI/5DT7iSkHxoVWyUZJJMW
UQY1aZkEyMpYDC1AYOnMkASRoBpIsskDzysSgas0YFfZn2gwdYnnFsh9PzgBnFi70T01AYqu4FiA
G+w6rhg1iYsNsBhrqX188kin8ysd1Y6La/yGtYxVlmBgNRLuEL5PBhPtGYi6A+4geClTVUNoZqj3
I5BN4/7IrxAGCNGNjPgNpnezDrEz7eB96Idg5iiPwi2yPwg56bta63b2fLDPIM6gX8wRD++R9s7R
pMnQkYy/q9N2Xbt2l5ooGHCqSDznPyedW/X4YZHaofEz080xiLtJjbd+z49sCUPVOnrEnTtsC+AG
Zi0YkDBhubdSsqiUTV41fL1OYPzrdZQYngtHlDP19mkWQpm9Cir5c0Onep6QUO4EatOCNDL43ylL
cZvxe+qUGZIny2R5M3gofDs59/JvguItfYM2gja+LvpnT/a1xD+5ZpFRk4Di8thmdxdqm22PgPxT
IgHbL50Zc7y3xFKKNyNXm1I0myEDM7wC2alJdpP4EhmjloEXoGbBjSeO7qVn99VcPhHckNhh7Goh
2x5UNfd1LxWZyYwrsMZnBs9MmGr3yoddTZa/ItnLFk5mJcysjVehRYalTMcoCt85K+kkn7FQI7mj
GZAnqD5nBuHefhyKEsLLc+bkfaXrVWEHV7VyMS19xd8UUM/mskFhNw/Qe//dlyS/aOcKFOmUpJ80
gJiiRBtFzTU3kkUj6I4abyExScCcDdVju29EondEk6BjsO0QuYREWeP1F25Id5NDzb+Bexv03Xei
uWkqoAfnswmGWbTEs/FSDIc2v5c/lhphoWS0oqNOWwNWBGW2V40Y+rht8KNa7uBrM5jsdiaPdQvL
jyku+pythiR67SpYcqJG7URHXFGkmlJHpeQ0ZccTbWure/gKLESk7P78TluKd9R7MZtRzRzoBxd9
PUjUnyDgpU6qyXMfipMnXlqhCbxICiuyouf8dNFIHQS2lSNUiAmPTuWQsxhzUGZ51ZqeFIKcqiii
DMEHzvvWO+FmtVVxcDnHPhLV5cwk5TvRmgCroXJ94SREoHZXdfUNiIFUMtVexkI6x989cCRe89Ln
MxvgmunPQEJzKnqjLD35tiQ6x8sDkSF3307qJD840psC8XREqdbPsj3FTZy+M+t7PEntUeohFWaL
GOgRdYKpimyUv6yR/YdoR9jktL7ajYzQwpIx4CJ9asYUhqNiW0Rq9d8n3vzW2yRE8dQdy45fR60X
WDeJolFtzLKuLy6+ZmJ/HS2vFpYI9yzG//xce7dmuU06d6mfi/dDDBd2Hw+NKDEKxU7eO5/DcQMI
yxAg/zR4ZN9lll2zx7NBHurvKOhcY28J/w6ra8pyV8ADT6hinIlwtb7wqcnLLZpii02i5J1f6zi2
46QuTtbWj0QoxhwcoEY+mTX34pyAcASG6K8aTJodFshk+JdOIeo1fcXegbyW3TDkB08CidGEPmiw
ObmJs529phEivuanXJJBf4c/mQ4doBaBjBUSnzeDqcUnLkvE/jvAsKBL7YkMlvHk4p3fuW41nk7Z
9B6ATBJk07mD2U12VBPrTmWyv8NFGXGkBBiCdOaVOIVJP/cBREoPqI7uvCmpqL4lrHwSFyhsLkd9
AErba6gvzStEnhYWlrASypmJHfoi+Etyo42+frFNOMsaZrBugyZ2+zvZlI3Z6yW9alH+iJW2YVKk
usKQI0Ny2KtA9YbP7XF67rpMLMOJvJL1ZQKJ4mffalYm2l4Uzi5Dt0vVqXjeio53ahnk+at2IQpL
mBY42rjxR82qJ2jx8FtG548kTaBbhNayh/q6Qu0V42kBYZAXGKrad+YTSy7kSLHgr1cNXI2izm24
XmjvUgXePIfO6Paa6JleE9jdD3l8q5GWD89BnZ21N+ZtggMisty1L8TQT91HJmtw3JiQrjbm6Brj
XcAYjSAvCkmf2v0x/DKAeTyAL8dd5/RSiS7+hFFiHHNWwMgmdgElvR73Rb+sGb8iXQeNbIxV42WN
XA3IIDqC/JFNHTWauS+DT8eV3ekN+YBQaGG2UYDoF8WqZ6CG1ePQ3cqSzO017V8Rh02w51XHHkbb
SoGuHw6xWXr0W+DnC/EDS/T5uYr1kzNuoUz9sHdupOL/E9SHanUHD6W6AY/UdOzeUPgLqQaZaRIF
FaW96lvDnA2iyYjYaGFJRDmqBc4P50fe7TF480w9nHVTyaQNv/2azTYgCZuSaya3NK7O+8mj76Qh
bixX1myz2qoqewqDBLVNGAmb1Y2YrdGNmOqJMlI7+HlFBSI4Rmi1k1/o0UKYCZ+m1IRwgPe6nirN
0LPxsSpAI8hZ6NMPhc3OSXS8aL6vi6H8RRmQHF+5u0E28fhKjetYaOTEqpxCOqdV6jJPlsy6HZns
a3TQ8HmLK0YGZ0ySnz9b1iN1MM3g/pauSL1YJAuP+gTbO1v3nDWy5joy+9+uz3fuVnKzudsjL6Ar
PVSpuY9EyE1Y2q0aW+tKGHFI+8UBl9oDmU+0UWGZZU0J0PGSDSy4pXNpWFevfU3RE7Drdz5VQe+O
pqHw1tm11JaFR38evI6f9+0/BBQasRKoPkQ6V0L7e7bSqpKuLWhf7XU5jDL6mukUViEjK6R4+thU
B2sK4AEjj1AAW3rgiQgJD52iPvswxMt7khIwDv6jC9ySe1AN3T6vmi1CvYpP6kaVtDFHSTW6lfRz
fugAmcMHM444U88WH1XIui1YqjT4zYVN6ANAmm7eXxbKeOXKeurD9mFBzwlP8SXw2/F7vOING3ld
imcOLSWCNnBSLQKZxgriCmPnbIoYuY67X6FWcVHhPnFp3BItT7Zlvf7/tlaqJbk38vJdOkMsd3bk
HmS+a8UBpkz7SQJMflkbwtSOs4mZNT2mW5FWWFwshI2Kz/Qof8fCcrERneL1p7B3OId7GRDxGBmO
6mEh+SyDG+mBNaLVPRlfso6656v9Ns2MqBlmqZBYwbj/neyovPsiS5Vul8eCERPGquByDejX+dta
VcNUJhwyUmmmHw0wQPpqXUGVkm4vyRJ7EeXyf5alVa87M7rHBo37OyeY99dFI2P3QEiykQTa04Ws
6wF/61n0I5WSp6ERBXm8LoRUIrysCNfd+zg6MSXLX8bzFh2p7s5mXBBQt3YEMkf+UE52IER7Av71
0gP/t5AEwIWiAQgZPfbtLz4/u7JaGyU4FQTYRBErZdMthgJX0S4uSFpRmQsuZnpxxOlIh1kILbQk
/qFnovM648LGdihHJ12YiO9CL9jzlpfCpj2G27dz+x0RkOG/MhlK3Bipw3P2SPF1+7WSEW9cA2MA
NFVJRUPpqlWYvNHGFFWLo2NQ7FTluiU8fpACZ724QncqYP1kyzSNpVakKwRAfWS3PMaEv/OvTf4v
bJ68ufdtDPR2yyzt6xVm5lhd8Pw7n+sX2kESAdvXcVoaiLdy1gMhj4aFU8SnQrPa8GG+eQ0o7Vt9
A63VDabPLnwccx4yDjEtyXj5SQOJyLR0sWfPQMxubGjStYWp5OCYoznOPvx7+Stn94zPYYy0mstL
E5hAsZw7Hay78HSdpzGTA+EHbVVqyKymqsLDtgBcN0yUbn9R9qDjRtG4XShZD0W00HngHn2ouaNW
C6dVYQzA2cWV8FYrlIyMsTQFuv8t7byea4h3YKNiZAci6RX4rj3LJYlWXNnirlYu9sK9j7O/8aT5
RKQ3Du8ioGbT2jw2a3jfcM1TE3VJDG8OEDtcFlYVVx5vTL/JtEqDxI/6g3WXwl/RaksooPwSBSHK
mAcugy3Cnd1pRxAwpw8cUXd8GX0G/oy4TWtzNzglm80p0C5V1aKapYtufDVojKjogWaYQAf8etcT
2a9STqjg1N9Bp4XoaWevCVfp+JfVFa+WwTTy4zqTlnCvsh6/zjQWNcPEzH1sEmsHlm/57/cwZ8zl
/rsFOxsDlF+qFPmsw6CB3ccNKa2v/pygY4yRWX/DOxrOgiM9liuVQeFst1qTkz174glvDjQ2u+qb
MC0HaE+YOxVREmBbIYxehGAOQgwkAnyTjKWxchmu6NhkTOouvgzyvCDiOLLs0w5GBrTtUeqek8Co
czb/xVrcZ5p3+/60CG13K/JcMaD4pAb1vdWCnlvoHqHEBh0Gm561jFtCVLN1/Z75RhkxoqmcWCz1
cDdwIlc4Y2BKgACCjYtVn24q40G7AKlV4yRK+iOUBPuGUzly0uRafqA6T1fkFTV0IcT/y62L50rQ
ze+C1iiODarEno1HqrLYdHm64U5gsTUpTfIwABQrBgr98Bg/yiTOmTc4CVbLV0NGiUPfQ0VtD6KE
bI/Hk//srbUGwPaCAipXvkVJHcadQsBKsVUJdFPJaVLKIB5iQkj9S3SJjs70ver92GlGtUkVJ4UA
HLSFi9Bcdrfd7ex2HclJ8ceBGh578fw1HUB3iENNAQojtVa+2HLEix/jRAPYA+h8f5J+lSYE7SQ9
dQjMtmyen6spb5MfsmgMt128iGC72ZFMThFQInTTNo7zTSazt6ryNrfNxPbeIm2DPP9tF4f4ZizJ
dvQqiLX2jgUmNYwru5/W4Ml4wrxX3knBfp9oAnRHEu31xgrZ9inXk3xcdp43hETVsENHTHqEj8w4
RGEXjiWOvcxMm2pcbSgbOy4QHsjLKfnMRIgyVo3D4k1+70wFuqlQGdFZ8HgqDuewN5cTWd90LE/w
tkZX3PlJY0CNpspZ/3GJ56jeKEhmHgylrj1eQg/YV2hbuVYdOCC3wb1bZUtkT71YxTlhmlMtSXTn
msjVijn7csB63MoA0Mb8FCA+COXD1QuWFkHHGiKZkAJovCwdfX7f2530h4eY4FhVJBV2Os5xlDi0
HIXgNxr52D/Xks/3TGO1KqrH23pAY/ZYKHFU0rzfWlGypBJHg32FAIBug8NEaH+thhVyvzgCzBYE
mmCJ11WiYIwFzaUR5oXtC7EzobVrlMFxxWZnxh1HH6cl8huDFc+0dAKi5JMW15JMd5v10WOOSv8r
lAgh1oXwOY2G8Mv3BXhN+WarizsYnLPNjBL1uqlrEwzGbinuWbuKBvFjFARpOS4wWzD3KoMyPq4M
3uYlmUKCkN303vzPTDo8CPakoaYj6TdyZEna+vZAllUBj/MSKwQlbbLYPR+ZdqhdA1/+Et9W6G5P
d29ZtQ8lsY7zSp443amgYVo4os0vk6nact2dicUd6PWqlJizH9lRZOW/w4REOdDJlEIG+mbnlSGi
qF7muMd7Y0gLwXlzn4ZCjSYkv01X0fL3cK3ZJzQruFTgZIhEfnvR/4VDwwX+7E9QtTtkY09tMQCS
Q/JC3kW1jVKQjHtPBV1L0umnJc0BXJeFYXgHPj361ad8bzy08IqJuvrES85ssfJFrbC2f7gxdcTW
Pgox+fyogoHV6DoEgLxLdMJuvJe+3RpKESUr5P5SEC2B1M0RnjuWUyb46psQCz5/UNXBXkHm+M88
GK+cQ2LGgqwZNXSutY3c6tDJA86UnBXzv/r2aMOC2R25DYT54wG6VXEOw0w2/xe+t5WOVc6WKV0M
AC6POrsztwkZ0nXmE3EioRocgUqzAd9GZ3M/ndWeGl8J8baRFFSYX7C8pB6cimIsyAeuS76SyAyB
CVuDt7EoQzE73W2AQEmeAj8xhiIIPfVQSb+Uslk4wRop8Vb0hJWjrtq3lrnMF7o6S0/OdoJr454v
GrgE02U9r9oRfRtxxEeSVEe4iOZSHaMWtHh7McPojhrne0jz1/PAp3Y37CVRj5AXMr5A/tyPApx0
XkBAhe1USOc/hLQLl0XNAmuFdBAz1V1a/1UXnQxY4PyDAmmc76kVyxe2YXLuWssOxo5EoIQUwadf
nE8ZNah/kGSJS0aCTrN3Gn2ESG0bdrNLswSCwwwNYMNtjpDpFSlqn/u+ScATtF3d+MSeo+GEP8IX
GJsCAvOWV8cQ/kMWT6atY/unBFQIMuweKzhyp67Z8k0lbpCUDBIE5wprgTq6CcET0g174M/+sSNR
BcxrXBq5v7CUSMCHV/VCdKQygFEhvIJBYczw2khO4bd22xzltAsCYqiyuKCOTxVYClJT60Mrx1Uh
gb84nGYgKu/nfO7/MJIwu2j+51XPgsaO2qKA1R47fF13YYo3NevMSE/glpwMmW2bhwzggJi213vw
/6ciEH/Wqd6wbxkjg1yekQ21guzNc3qGGZrzCmEU0P4sLxX22hpfv3MzeonrwAz8FUGoJEvtSrPh
ROXF+p2LB7TcTquP1Kj5ASgg9lgCmN9A2U6Hypld7/D2FAzBSZd2k+IzH+jUn+2b7RE/dRj/USTI
5YnQ0l9thQwwGKUpQw3KIyBu7l+bzNRPwhQraVku2xkhw8oKCUlsQ/0ghIHPjfKkT4sutScYKQXr
pcWqTAc+7UfPOLAaQHgaNz99pEHyrtJjhDjaVVgRyBO+p3d7XVgQUYE3rsorxBTxYvmWMeS/vlRC
iJFx6iviYaJk+Anv9DMsYhUpNI3zoC7VtHODeBuUUhNS0WCQ6nVdoJvyVGcYB/xVEREBoM+6rtRS
oGM6FpD1e34EVSXF2z4m9cN2UeIPV1vJuTrRhzpsTGExW/J1Vn/ay+MC3cozMA0TpKJvtAST64Xy
w6myXlu1GmIRwZNuvpKw0DVvHGw4flLNJ3OvtgQD9hW/b/RxVqdgpMCuhij751JsLfYR1GavEsGc
Ka1Ma71H4FoBpfomx+s94JSJJejiNmjR2ut39yORjm0XS7sBri8issUUUjqEYExd64vH96OmQIEP
3iHWiQEHLwTrg8kYrS94nYn9N8xqd+Eu3S+/BhITM6xwYYv72HDe55MIhttFM74X/bEKgSjXbhq1
LYzmUpT+SH5Egy6dzZdhswBXuUKFM/dWhE4iN+5bwcqnu5v88425mrWQooMY0FVW1bXOS8u+v4qZ
XXhch6AfqSMGz4C9XXbLI/jwfLC/jutsinBXcr0gcW+MvxGKvhBIoLpzlE42aNm+BKwZt+C3xFmQ
k4yLmOtPLmBc3IoRVIKy1a/Hl016AHSi/QpPN2MqcowGWKcTxvNJ5NWdm0rRDL//aXv73691Z9KY
lYhmLcF7G/7BHM4Ngz84gsNUYvnWURZaro8I2EncSAjwaLk0rqkljKxa2mg7+XkJ/31ZzrPKCCbP
kOzpKKRIMsoZMwUfJFkccKBgJl4l2yL+DTLPAoyFSnoxP+tUt6VY63hkk7K23U56h9tWnj0Bqtch
qGasydp4VI5ktFn/r1QeArJ6PDH8y1aIpR74mfA7Polwi0xbQ9MWun+XEu37dnrcNBS+DhDFS9A+
F0OrMdv2RiKUyeS0hpi7EgjpZ3BiKQUWg9eeQ9T9jmDLJJjXKweQiTDy50xJ2CqTKZaOJZNG/Akj
Gjtz9wUUTnOgz+OGLjRNuHBXSu3VnqZogIXhRb87AsXgi+x51RPxND2RFHr55ln31Auu97z15OwZ
lgqa5jPw9jAOW1DyaFL6XwTo/PjmD1mVDAqk2ovrPt8ZOWWY8Awyodwlypt2uFSSvJYLf/LMtxiV
L+q7RzG6GbZYPJQvl39KUqYo2Ie0dJ2NoPY8kyA4vRYjHfUCaQ15inMcrGEbbjtrz2bNKYlXLVxT
MNA9EJWzplmLzjlPbJboSOiORliuWTjJ4pm8Mq+ZYTOHt6MACcCHry9cUo6q8iovv7lZJQYPBWXx
/eAsCxmQCfWg1pbNuNfiHgGF/3ibWTPwUEwK1QgPVn94qUslFt/tye0TW9NlEWOELFVizmkhqVFv
lxRy7DY9d00jb6j7bqWSgxYOUomQz+VFhyw7TJAneMOZ/32x/kwZWIsVM63pNcaMR6DI80JS2mRX
L9FV5O2CtdbLpnD5SGIMgQjQmlrlQak2z77WKTsdZGMTBKSbXlZuQbLgbMFTm7k81SMJdwRbUfJF
IJ43IpyYs7XN8vZ8tnVXkuwzydMm+wNEcpUk8woOS5zsN6Q8OZyaKsegPANXRd//a4nGsdEvJT1A
yV3hW/www0GnTPCpQouvWIGw6uoRw1d2szDGl71JNmo6e8ip1HiCFTQD5HgMyCe8JG7MK3Dk5/E4
4urzmsNejN7vvIVs13mhqVp2j+U4++85JDOy3q1ECE0M4VNjxPxEvuvqN7dFPKNvCsWio9pdJrB0
99JEHog+NQfLoIb7qNsUafgvBw+acaP4CUdGi6abUwjj8hzpyO1oVrJl/oGJa5LU24CTNPAdB8cc
1UqXo1zOEa5hkGJ/+xXfRePHfN62QjcsMIOPMvgwcYUt2qaVl8bNYRFIgqNelartJHIkQZ9KbRny
I1oWUdycRU+H/uAZWk0NQdVK1IMyG4yLGoA9DWii1BbMktjugf6n+qcmLeMCCNSYR2C79J7i0ne9
CGR45l+iYqGl+mt/R17DJbwWOrClZ91xNqrcSuMQ8rJ0T7dXuPLXCzkKzjxzDYPxUmNlw2/R2UqE
tWZDb/5gsh37IDqCsSPCjNFC2PLOUWzt443JqrUvEh5spxwQoLJqBn7XBUcUvwlXsLYqcUQAnTk1
vNHxqPQDL+q5DNTJW9RNdDgwe/biqow194BdZXNJDVzyxgu1wa85amfNbs9iKxDWbfD3bSltqwUw
ZHRoPxUAK9vy/S9OCpcG0S8nyiJWWh+l7t5FCj8VcA9/ItPMQuiGDBuSrm3ZxHjtCRZZENme0S1/
YCdIpRXUMfWyVCMyPxflW15+chkem+Y9nSpId1soBPKyVFV7Mr+cNCSxNjxnCm2CORVGc67Exlq0
TQyFFDQYlNYliPBy4A0SPWC4uOQuObT8QMNBWCugDqgjsFXBFpZvWCzhBtvltrTUINhDGmkJ4+JH
93K2TQ7C9rzMjIzip82PZbjGD5P1trxewGk/0jc54i4aebLiiBMkw8yz9RwX0PIHYT0C+b7Xrral
+LFH7n8LvbkwHR7XHomdfZxPdeACBxy6AalRE65hh483tTonot3wXNyfIcjwUW2kVVjR+vNFmCt2
ug7DU7VHjj8+f7WNPe0nwWsjgUqNFiO9RUulryDZ/ydJwPiF5iSImOD8wUMvUUZKb+eKanhMGZX2
DgUXIdCO2d7+tdHdooaCEqmRlQKsYqKp9UB1D2j1RRm9G6+R35FlRvbpKUXOA4MXQxnH6e0QBZI7
Z/ASHk+ERK6P2/yNa7hiQlyGfMzSMdmjDeD1LEYxq7JzOTN6EhUlB1G7ybMvpYqBhPimCLpNPyoU
6kmuMbKwehVnFIwwtNLeE64OyWwcM4gIir0pTd4Ez8Xo75SnYpaIZgtcyyZDwRxoxzz0MwcN+r2R
GscKU2cXbZMPfiAxB3J34TC+5kFaTZ8sg+BHmZygzK+a6aF1zNB+GjxDzgZv3AWUuM/RQFWZOF/d
zYD1tnPnUm8qEgmn/1n61XWSaVx6OrUnYrmAnHoUXdRblwvcZELwjGjOrfawAyRU3k3wXZk1J+lI
V3eVnCaZ09Pw98YdBD5gcDCjJQ3XYFtxjhwJj9nkHXVYmIz+DDIBT9jRRkbr68/dkPN9qiQHqs7L
UEQ9B85HBy0rm6MS/g2MYnKHbrcKYWIOTe+7ajdxNvW4MwWsUlQbj/x5PzSXHj2pgbjlwIjKIKEQ
RMUCACsnTMPPtr670wgLXMtLOs2z7rRvfJsQ9z5aOv/4PVeLhMn/NfRgaWp6JxOZHNg5y4aZBXP0
fupRMnsApcbrmg+yWdFKFKCRcLU7n7czI+jGDybaQYWvw0WuU31+Qre4QRnWzgqndUqarTKjWfmO
AF7vrtfx1nFpkR9imiKBhjx0UGFGoDJb4gIWczf+ll5IbF74Rhym0hjr6AWeYBJ6wPpJe+jO2i2P
FDBT6o5zmHw28Ygahaf8LcIKE+tLd3WVpuLiFm/QQ4WXM8QUlkpqbopvqyxjbfyuZMLDX3X8Uy+L
bDYAfl3QS1jb+OwbyFz0Hqqfm0zLRFZyqAKo3w4qWYttR1eKHZLPG+TqC/oCH6ZKUYzhGmKNOZwv
U4aquIa9uoZpP3/PkP7QnSPJ/5VO3SBHx4MmTXElFdG4nb2z6amhNSQvLZaCYHIk/upCoJCVooSW
YToneGt5jCFzBZgLAhcNRq4hcdFxJJK85GNRSPWrEEwWQ8rpMY2V8o+7CYn7gVLriu2xO4KQ0VZf
QbD/dng7lrcUaqiGPLkyLDEnjZa4hhufknJWbyyLhfwUtyuQNJjGBG4YvD8HHdDLpU4p3OJxPPL8
uXShadJGr9yme4enFxoHjtWwpxUJ85zN3GaPbHJzM+gLgkvo1uViuTJh/hoflo6U4aUJc+h+miii
r+tdrvc+ZvCdf9mAmYrCXBF12lHyzGc+bGFtb0IXHaOJosA6NKJHhjKh8jKAX/DbXwt94XJFHLhg
U/4tnOfYGCgxklkHUeo1XC65qzL00OV9+lxo+NGjYpMc4ke5sXnKbCK/JfQrBU7OcO9lQx3F370B
gAoCrCa5wK8tfvX80VRmdPjzJ3kzH255a2hup4iinMsESsM0U3XWb3KC2fVvgKnlSBGpXgQi6RgS
rmTPRMUXzB0Cy/V2t8SKEPNRCYyP9sSu2jISwexDbMnkOxtNtX0O6bdDO4aaF59K0paQ9p7Hef7+
xxl98gI6JI0xQapL8shkivmcLgXdAXKRCppgPuPlJ3NUltIzGLbKZ8gTAJ6plgsN6DnPOvWhWIax
HLiiLZj/Egn29yCcUwy8ddv08TgepiYtDv4hOGvb1lpGDimtR6EV/rlmAvOXIE5OOBDQLKiCbyjD
kT1xy7lW/x6TsXkRlw/DjR/W3WEv6H8j9hLCkfrOC4JyHf1q8P1HRNTLv6LR+/0wQC0DoS5RaEE7
lLzNDgZVyM+N7pn5lFX1fsRJu5CRZqmf6mDQlFg/QidGCak+CFEO1BbdcJTX9BsdzAGvsm1k5TqK
IBGGVpoc+B3TCqcYeN3qHB2Q8KzaYyK7rP1AOFiE/IftRgigtnqecXmnZXTsxEUI50S8F1Y8PqlJ
7uPM34LcQeGsk4HG38/cjdbV1qdAjGz22JUmKMBXKL34V895ylhuguDLcFVRHjGnLatgLczf83pg
98mjgL1dvXSLKACoceJExJkQRyk3ylS7i6obniT+nLFre+9s5B3HZftm8wHScGMt3kARPyl+yNJo
tDv2DryGpAkBExa9u2RZPE9lUQeOCBKs9Xq4BZl1dOEwManh+jthxlNN9nNjfjN3w4uVzR1E6Ckd
5Rf+x+IXUAGou82/gIYxCYMP384R0U2uI6r3nwsIQwNMsEyHUU8lZS0k1zMo5M9r6YoOlf364DFv
PhEILBbtuyoW1RlXpFUpxuJNAcuO9BhDCcFjadPnK8T8YZrBAsisOeQXDDKqcwGkHO2pe1KIy2pL
RCfeD5kn39GyEZxR46mCPS2Tkf8z7uEIi8sMCLocAQZD4fLsiIfmkmLu0p2SoXf5bOTxXUxlY4fh
KDr9Hx7581emE0JtJ25PV4xgGtfbvNhA1krf6wETkBw9hg/mrjJhW7se68mWTMTORF/RWkBlhOwQ
1fdB168p3Eov8XZL7nU9nahoeU5lPCW/062GA9OwLx16pBgwN61JXBxgWMQCc38Z+35sIWqSi6RB
MZgGFtb/ZzAoWWFThT3e+34+sUpJoJ5GVev9maaMJlc7f0cB/+TG1rigwZn4X8T/UMCgjfg9jcSf
TvL4H6NkjVeeo3atQIaUzN8otNpIe9pGxOdJ+1/39HQ0nwTLRBXbLvfnkFwqtKFga+PXcwg6cLn8
WCM2zsdcBiMw5GTiUQSUzXQoOLmTe3KEWMvD4swDnqWa7lNVhU8fb3VVBgpZoF+C/KQe9bhPSWqA
it0+gIDjKHj4cC/Krdb8MzGhgnmdNfO9ReqfUFtROEW/le7iqr6Q7QfiCrqzJDvB6EILgjkoL/JV
mAx5ykKBkxoxI2tb5nrD4e03PypxV5J0NeqgS+y7deQqk8VQbMihxVhmBNKRhniyCWdaWbb5Gn+i
1mDZed/EDKQu/bZQUBH9RWv4vc887Bh1gJ46FUaUTeEKnHCBowBDGmh+BmF2snbK1RWQJ9EKfG86
EH50KA7/5AHCob7qR5Oe3/5CT1ZzAnGrmju6DYLzEexVO+KrZoBLN2dskx1hZfliT9LvGoJmmW02
KfUxM7pbtK83+keb5Un73/38psCPLvezuEWFmb6vf2Ld+90PuWhnjaPGdIMgCVSo87UpJS5rxNhb
rXRMAFLB8h2c/HODogvLHGusj5RyeGZOEeM8YAMcH0hwYzCb386bvwsqY6MQzPXmNDVhZzAJ1bof
gqH8chuddP1afptUiaoCi4fJWnV75NSFAi9D14st4GjMVBZztnulJkH4qGe3VQGmc2A/bIyDiRk1
BEdoC46Tw4qsQJaU6wBdTLfG03hqN1IcQXuZcbiMmrTJ/OOfDw3hpU2ds0b8VlbYKfxhVvhfZRzk
YD/me9sPb+7x1QMxOXbdSWnfgmB7L0WAWMZN/lRh1kiuTHj2MjKcgX6+IPCHI1WygiLHLFkOnRdm
/S0QpzK3E+9iucmgcEFdSbMx9SG7Y+Y4zIAyzJfb02yX7KlKnlu1bVhDoJOrWbvWtDvkSV6osL6u
/Lh0Uw9m/aX2K6BH4IrPbWyrPrLaxx/2Yv0PBt6VtJtlpDikKYc0yGYgX6VRd8Wrk1tgDsFCy3FK
SX642lH6cauBYO87sIoQ5jYnOBvCDmAXkq7y6r0T1Aa67tdygb0ZXliCfqCUJRV9/lwLVfT9KHIx
zfMKuDWTekbXTUi5uNbbVv0XYW32xbhz81FgpF406g6Xp+R8hFojQI3MU/lmsuI2BMGH/Go8jK4p
Wr+nJ6urjoyGXnKZCs3gvV/iOjeDK2pgIJ4NqrezQkvMhijM+Tt5TIt30UuQOIhk61UoB/YZjVFN
gq541Lr7klz7xXu42iVFlvfL4DFuckWKS8m1XCOp+4htVbkU/1LfMziELb4p/H9VDalzduO9geFl
qHTpgs5rlWc7iVS4LMrvGh31Ha+u1mCuMVnHPiP9Q2LRmx9Mb9LAMPYfgmJIWJStbE/bFYCO4ZOl
RdxrtkoMiCx0MMdKNfQsnIWXwR2gbIs7575IVvvqhoysyD+E7uXoBUwmA/fKWV0MUNJXwRkGJbdz
xt6XvxwLan/Tjlckt5FJEORg7BloscOQSzL9uKuFn26j8jh2gbt0SJiBRa+rzpcp91g/Z7OtuRYY
hSqEac98ColTFjZb6ijt7DTWrefO4+4c/bzmJ9rO6IA/QA9vjS2wRzOSGRZDryxDr8G2L5VZibXr
tev5Hzx7Nd/us0DBE+y0I1e0NDX0nIJ5/Z8RqYJV/6azneEFHfYGNa6Ov9I7LSiZ6HZHsUkriGau
g6hupKHrexnwAXCods2DFpfEiKFvxLXj70lyt7f3SWt24nvYaRMyYJqjrgNPC3QszyPk9ZNwqV70
t5JdEwtL9mJCuqIvMzvoJcQazULb6QDFrlkvp2rXIssY2dtrZ1UbR3PpW4oKpoPii7FOJ4YJPKkt
8HUzNIRzI4Ak+tHyVBAuouB31vdzoqGaQVQsNkxfbfe84UdVB0nWeJ5dtgju5ZXmau7M+SrZziYZ
hyxN2EWFEzcVyqAdMUrypiXIkLhhTwZ5MdrVg+V5/N6xD9YLS6KJ7Oo3b0DwJt00k/B0YgT7Wp1s
od2bM/4Ql5xXTu0n97/jmSOrHvVq3Z7Dlk7cPrdjKsGsimCfP5yoEy+M/pTyfk6dj0jFd4bW1XuA
bVhJxHhPk7EZj35+WvKQeP5xnZbx/m/CXPhHEx2/z2dp68J8ImD/2jruCpg2gzL8qB0LkOP7+twO
9YivOZNx01hi/BFcgazB9jT+kLDGl8ZmffhsBT4HsuqBHH+OgrioWMqYYq6cazgENVjWqLi2x/eZ
UQywE+RFdQc0Q4A+NrM+WsI1JNlVZNbmXljTn/06Gnw5WmMK4hH9Mg4tSlfvBLX4OX1Da56E+Hh7
SpBEHaGxMmEniH6f3PJp7JjnMtL1XomQ+83hftlE6v5VaNVFECJEs/UN0wUXQIrhmnUs+XL3MiUX
T0VHMMgzlLkyC5zdjmFM1kYwDNZx2kPkEWGD5ubD2PV2moyhJ3ZC2qKRdzq7RpErMu5m+ojBuIEo
EHnam0baHwkyqvHDDR2HHNP0dbAiY0k6Hu2doGxJ0KH3yRsNX6gPJVYLesNLXc+QD7BZO7DFq5AE
fp2jpywW7vr0+A+dXZy+3TtRk+R3Fl23hYV/NJyfv/1flCeTJxj54iN19cLrxIPNtCHZT17bYuUg
bMmOk+q21R9P3UR/pxSW9xu6FFbJCmRKXvicudF+UbtU/H9nFycr2MIuiMdIiii/hg2B9Wj9qFTs
sSaxBfANPQWiCon+Nc8of4mXWxt3LdI1wl/aZnrWZb6QU+iyUgTzi3FueCGg/+pWMmNKrVCpPH9z
b7o5oiVCj/f/CnxXf1edDEleHVLGR04gVVLLRN7pHMnxZ6I15++wjKrIcrCYzyPkPNkDWMx96f/h
EiEAeVp2WNa5P7oz8Uo9+XygZ18/jzj1fR9rBBXjA4fu5toBWb9JMHzeHwzK50dFm7P5ZX0t5DEX
4XNq6pXmOEIVG3MMge5ViZhYuJ7HN/WcY3Pkbl/y6p4CYp296KeZ63LyYD251Q/K3In7ToZAj6nL
GjqfGAFZ6zFpwNiulKuMiko2DVwV37aOmIVhE+8VgOETrIcWKmgTvU6LoLWJB8ulPVetEGIjcyNh
bhKAQepPwllE0i3iiN787wqWgE9+mOqu/Gh8azYk1gkS5e5LIto8w+1SjZvhdU6xaPmZoOYsXh7C
+UMl39dX1m1I/BbqE92qG5TOIv80+IYJzCSWvnS89oyFQYqD7h+L4SMCdPSp8KO+cEUJcP2RLQkx
DiwOrEx12p241rDxW6xmujvGbjfV+SnS8bWTVOnfIZvC3ZTbfUJGCUjb96TbCoU6hf9ByGXaJ26w
LJENqi5X0zmqhth71dcUNOJn1Rm79vC38YzIW7CZgNf4ne+0DmdISDwRJH/cqS3Y1YZR8wAL+oGA
0Q6DS+WpCn5wfYJ9zfXe8UEbl0wnEWgL2KPAP9SGc28boRrQSbNcD4NhIPuvbfa2fAW8ioQKtQb0
tIny1zS5U+DCM+pgt0DFRT4iHQUQDg94AGFk79MhZs1A7AGHHsF5IXFgg6Y6IbGtfggLPZBiikf5
HSOD9weLRmbEy8IYXsji5aE87Rm/RprTURFk3BHPf39/bIiyr7FoxfBzv0JZ3YQww3xfaK4rxkzq
/KSW1yKKulJ+chPnZ1Peyu19Bmr+veNHPV3msYnWvZjwDhfStNwKEAgcw7khvWzpZQQth27OBtye
0lPUVTPUCu1/GHmt1QhUSV7qGCf6MqrypUhdozG5dJg7S+N7bt+AzLa1cT534kB4PJIlEAO346Ux
zbgr78UxbbiT8/Z17Zwmhof8dIXqWEqBWX961sOLRm65w96lWadqjrenbW6izvlpa4hlkpeF7E2l
3dRDh3NmNbkra1HRGkgLEEcDZaprIAMZXsf5FNQ/aFN7b/wGFT2YgHYgwC2jQO3QOSN/S0Kyhc2g
Mj+L9RSXUDXhEH9ohAw0xhXgan8v/IAIlFQZHHNSDvuMP9pRrRD1eY9tRNl1lNWpFnOagkT7Xi4l
yKZaEzvgNkdsGbTvAX/EXb6ZsO2Pd//BZKXA6Jmt2LO3eVF6s0AESetU/ut0XyjTHV6kZ4oD+0Yc
CjV7WXnZ7WiJPkiwDHmN1TAm8RsiEbZDryNqkfU1fUJ9Tnu2dM9ggWeWqSQ+gr78+EAhul/Sp92z
pdQTqERXg2IsGGzzGwjhuW8pYCdOskeSuEClpAM+VN/fhJUeK/8758/tbb4qj/xa1+wV5NGJAxiC
CavYFRqBVhIs5RSU8lOVCGqTRKz1au0Dq9hUg1xYzGGew/t/u7+/ALSwtrcHcCviknY0302/hLvh
VQA9UVDVG+duDvAz5HD66RyO8AsDXt4yjbGddvQ6eqnheyXSHlNjG5rSCZfoDN1uOvzZzxkI8mpk
1hmg8KDpq/hPzYuDBsUlGOqYCfkOcg6Dq65+HuPXYmITpaKA6c8R1xItcGbE1iDcjwR2YA/W6sGO
turwyzyjs5C7QgY7KF+dBcgfBfmQ/t0REnW/ZT9Es51jB5TlCenC3bv9mOKvYgcCRzM0vkaZe0lG
spCGM6rPky7SWwMQvlg+lpIXLm+3ZachzMB6TmDb2Np3R7ASKGaZ+jUKXlGkBusDiw3boEVFSK26
hHRFzPFczd3lSRhyhRISSEkBZQLCG44DDjce18I2P234lQT6Nue5j5l8jmVGAMtllho2/qe46drV
5pu6rNro0YwnyZjDeoF8Ex/7GI7K6B6+1t2qs11wFdWhNsjbDsINqytBIKWhi34tq+hR+l0/ixFh
DZbucyFiwFmk3A+nyGiREpwAzat/scpP772Jnzdeats3PVDjY1MRbwxlD3SJpJAogsaKsXLHhmtM
I+//TyaDA42TA6SfrAWEXF16WvNwR27QFX0RmdeVvzkBw6KyS+QlVkmxTCYa6o65UjlGB9Wk3d0J
UOhxVQsKMpk2JNwiqM6icfWEKkr4f4wxvlIO6Uk2XmsuDGMGAwuUWj8jJJ3OwIpfFUuiWrFFNMKq
IIJzbmknQwGwJ3ibIiVWgRRVv01GpmCkfKLrDcT0PRgFw7q8icss3uZnCfINwWLoI0HmRHx0F0ER
sVLgGPzHAjnNe3Ilw5RDZpemEol53dSCVL6c6k2qo8ySYPvxc2X6T0RxGV4wvuLZYZmbByG1N0E5
desDhb6PeSYV2YYtNRD/nukoQExiIKUobaH0sCRQGfSjpFG5iSaz9AFYk7SGO5WbxKFXIVd9IAsy
gKaeBF3iJVC7M2Lxuo78wB8qBK7KvLJW9GVP4ooyzQTzD9aaHDwI3Grrbub4fJAHI3XU04QF4tGG
V+OIgSXjII/GhwwIheAXkG9P4Q2aZkWQDf1HSJf+w769K7EHHQyxl8Lwl9olRr2j6liJk/F3YR1o
H1nl8p6ATOHI2sIszJu7M6lFCol7XRmjM4v8IoYE2qrWevYHd6jxC3tYvX1gJ2A/hQFEWNM4/LeN
H7/8ZR63xnRNFz/wwRoMVHH2G02+67chetvfv2qJJj4JlMN1yIJKpnulMu2V9mzDbMX/vhQrI6u9
JXLftjo5EpQmc5BMV0T/JqxwIly3Bubx0IN07cbLDVTsgYIC7AfcAp04pufmfFEo56S8BTRnfU6T
ARzCjriKkW55Jf25/t+cGIVfD/50cVDrM6szbTozO3Dfdfn0occxuQIUnNlYF4ah5+lGCdFK1txG
SXAwo47FCeoIxT9ef0Kv8GRlEtP2Qupnx1FWCRvKrVWQFsTcoedPmwL65ry3+ARhCtqATGiwjbao
gqinMncGButut6aKCwF5iZJlxpna/8KImnRviCAc679EZMAoOFKkNJ4NCsjwuVr1pmNzqAXuMHhm
b2kpLSNDBTzGLAq+SB5WugmJZ6VvkbHKPr4OqT1jaaYyVvgGN5+3OvMG+/WQ8vQCBWmYXaYygS+u
cFDQlHJ5EG7weGSyDciQt4ksaspTtMgtQrnNVGkKwtzEkNzUg5NA2L3Z28DiFh9IwrhmGrCaZZw/
D7OqM1/5VEwZfASI+WFDgSF6r1M8ul4q0vynTeX2Tdrp4NtIdjts+2qEheNjHGIGFE1VmjABnkbe
B/oDykSZ2Qi8qiVmmRILXFN8UhLF9GS9E4TYncXHEhE8pdVIrF6YbGtHvjyPKOyWI/LYg3bPEmeF
TnNcdmZKxn0Dsq/AoFv07+Y2PqpPnxcRHZgd3EyK2+2hktBD6cEKLbVgUxAVnF1s/KrehJU+uawE
byOV0cqCK73QTxmG7aNqae1C+JGELluqqvbvb9W7yE1lbOYNaZPxFqr14Cd1HdKoEObhrA41+puD
fnUdhOOfUYN1VO6FgAK7qkgHr67KRZQRRujjnlSddgWuVb0Us18cdTXy6cBaQ0DoHyPp+UzZV5aO
FJ1NvaktGx8nKMWLiQB4G7ZOWgviy3MRBMzf87VCtRORjsny4DLe+JECbmzL1D1NUl9gGc9WmMeg
7x68BzjzC/L1U3F5DAHh39nlurAi0xqnUbxauNgPQes1WX9FBsgZUHeex/NjZTKNx3KdJBmM1hJm
zZMTDN0fKZFpelPAsQNU1ME/PX5asUQBbt9x6KBjZfQe1W/0Q4MMft4Ff4Mf3AbB/43yk95cOmNo
PTSp4wThVbs14UiKz0VBI9asOScnMFvlAoji5zdWUZWaVcfC+OvLRs3jiQASpUFPQOIUBJmoCR77
b3yU0FY1bguZ0wRDcUrX9gGpArj5mkhcghet/Pecq5ocw95Ex7Q3inxbuymQ9UqSRWCjx7omLpZs
73PKQfR8TO3f0bQrXVHSM63A/9b7UIudHP8tpENirEvHVXOO4D/hFzyVzVwVHk8M5kgUkDnFsufO
lE5MrurwM6mcRnc+TBZLOihr2GOTvX3HFvs6yKJ3/8NkMqdYKhLR/50zi5dMxcxYWYGozp/s3H2N
UvrwcUtKw0mU++okRHyPeDS5sYibBM9kORas7kpM5KcsdEfAsH4cWaIQhTmjsv1wV3LDSydpmP46
KaadvNMcu6zclqZOYsi6JfdMPVvRzXkyr/dsK6MJsoM/szb+Aux9XQgk+Tpbj4rJ4kpDmgS/1TD6
RCMW61MoKLMF5NoBeG5NrjkXPxAwOXURf2YiXYdD7/BfJsjP3DtuCQp22VDzU1mlcakCwBLk/iKH
AvZVOX9PJgHpbCF9P9ZgziVn8S8l17iWJTmlFLqlDAXGUy5AfPCnExpkAGJdH4xhGigJCvoeXVb2
oS0wOXQb+sd5G6ewI+wlCGLDqBrra+ldhvD8i+hOHerI1iu0QzxXnso7XAdPYjktkywfQgO+kMOD
q3sNHjkxJvZNiQ5b46uBBjYRWhMJ6Fk2m/GSQE3gfvWHq+7wVpZxeQjzhcbNMWZo9IXi3CINM60U
byPf/TGOKy7IpYaY6UAF1Cvz4MMKfcomARNmcLiwOMXcg4PDS5O7HIWKs8z+2UbtGarpuNMoyZ/+
m03nMFYAgfpqeoBxdrjevfm9BpJvf7k+kWvNkF5nfIfacAzVlTi6DAAp75x9G4ufsGuGKBaTU63l
/0GgjdtxC81qFnBGROhQ7sPGXR1VdfhWZt774vpE1Wg2yjz6Dr9lkSoLnkBZaKUjGnJd+tLGRDK+
ip0dPnWMa53dMYbrH93ywOw+cedILOsrn83LA2uRVPL/2nUCYR0PR54RGoz/ItRMDgIlfqhpaOr0
ybKgVLkmMo3/w4YrpWodOvprmFiQP5Etczr7abhBfEQ3DMZ1fKdrr1NkhKl7jCRP//KEYIR55Zty
InL3Bbx4wdh/7AMbjYO1BhVvgl6Op9uMvHH2mjBo5sRjTo3MyNu521IDhBiNe6OjNIbQyQRASDNB
QmThSsy61uqYLiQ0ciLy6QqvnPnCbhr2VhMyJZ5giOxfFLVD14k5vAN6NgxOdE5ZJp7M3+Ia+Szy
WMMwCbAR2iTZ7eo4zqXvoM2UMpsC+xMgaijviTeH23BgVVDQcwUO8SEMRSrn6Md4A1PxXnTSYdpp
WUPePhVg5qPgz9KCnZAXzuabs3TRb+lCRMIHQ6huc0tmAZxXbEMs6Pjp1tqZAu8Yg8XLyxe2wfmy
FotyyhwC70pOp5tIwMfdjZ5tfWSzqXe0unOiwFcTQ1Ztq39Z3PoEZLgEKB/FjLQHdkdWyiCJ4KVq
yfgSv8XJacV8So9H7aZYiftbp2/9BsVvDW3pS2cw3b0xv/8iuYSF1payBybovdKgxKLbL7ukUqUR
FjWM9wlSvsq0wLipujWj5+VhBGR0WHhVTCM59N69crWAxLJSUaJbJ82NfX3tzsqhxVT8kpYDxaRF
SkIfMCiqdTpU+Fbl+JDmgmNo8r6kNpQP4AC7lsaxCDBBrBCPmsRwWr2H/z/qZeL9EACs3o0PFNXu
UkEjz1NCVuBpV3Ij5ehoBPuk5xmgVTyIbRPzo/tEjQmol4Ol4Vsy2HzH7cFpCTjRwJnb5P6s45Bs
VHefQl+/kXcTSOLIvppZ4gBn8nIqCWbE0K0ehCCsDTjSgXm4Xd9P0Jwp//bWFiyDkoADgbcOERi3
4q4bW18xE+l3MqsSVhy8aoVLchZLQx5rP2xxWeP5oEuawJ0DyR4ufAiSosewb3ixHx90Ak4f/7Lv
1s4XQIw4UFF/WrYgLFnC4RU8TCv9MphMKtHOxfj973DLVexHzKnVGHt5UvJxnESbAPa75hrG6p41
Ek05SDIO7U97GueEo00msd2Xb5hLxrB8dgtFMsDhaul7MmcQEfxgICbX14pi+qye5Ojivx0Lhioi
IuUsiszeCwSKuIpkN7hh/3tKJ//uvAXehyTHukPJOMWZm/qsDOxTwy8i17aMXySp6TUDiR0Ov2T5
ob9c6m6tpSCqk1PlVHc95/REzkYZ8mstj9udUHWycmljO7qHo6pNa6JSTlBtfzuVf1wr75eBjimL
Dee+xEA32eXravcTR1M5z4GtuHRKYIHbXLqhpOjvI9MaKG6aIErqLL2uwvi8a0Yp0fcWgapfyLsJ
sQHuWMiO+Dp8H0AIjYuhm2HoyURDjGYxr6mOsu+GBWuarVVLj/gx6DLcw9QbNAbgkgaCJ2/G1HP6
kI6y2TdEUvAGNY4j5AypVtuR7nHf3F2STv5H9bzTF6SU0+YosOrXuNL8NesuC9pE+R0VTxHlKFdT
8dQUDOvqN9SniEJxVBP/x7UeWUSHJfmzReKzci096X6t+KyabE76VVbnn01+tPy7GvKvJPTheSj1
Dpgun4JeoZ1PQ/NeMfWY9R+ZJvYyMG10rLChmdmvG9SpoppUI0xbEt2gNKxbYNwgLPwlMnpbqS9P
2ppGwk4la4GkcPw3Kor6DU02+aIHKEGa42xKP3hicUN7pWvAmPUXC0neNBYSn0+KAa8ytenoUuvW
CcwTdB78OwgVP4ONHQ5KzimB2iSvNGJIAXga8rUqO18MXSA2X3AxWUxRkKfEsaTpRtNde54Vdjda
twPTANG7DtaEVIBzT6bfDsEYosrNQnWoVu/VuSnBhIQYhQpxWa+2VGfuYtYsC0jrkVSwoMKGbnOO
VDLx4CGaOqSpSr2iqlztRhYR8Zi8EBJgLhCeiUAz4y7r9vFhFX21kn0R1B0eDii1JevtOQZSfDxZ
XjgFRdoYiGE9Sh3ZnEaWvvcofQ4mEEDxQrru/+Wj5jrqQPeq4TnpypT+Q1melcbc1nKeEzmC0IZx
1G2Ut7zH7J4hL6UpePERTuv6zDS2zGvvEEdJKMKOwbxElPqDDBRhuisbaPmXq/i/tfZMI8b8Toza
rP9i7d8lMKhA7GWwwpx4OloxuSlMvZUNReGFG8aMIipkUq3vXv2asu4KfG2pA0Mc6oKKcVxFhgCj
CNg8yNXGpzACOStvG8HpFJ+el25RExGXf0jrkDS3wgnjhtl+1zVvDZQyU+fLl4iu2QpF/6MXgUJA
nCGmEwdfZbdObuRQCIt1wq6eD3Xnraulps35KGGJxWab1VGR184EoQ3lOT28cmCE2ZeHqy72Rp0e
MNWjLL/x6Kc10YHQjp0+IvPcW9TDT9ckc5UK5XYDUEXpl5x7K1bf85iOVlkydRSMEGDhdA++ZYHP
WrLFFDNNTFA/XOGT868RPr6bhfaOTWSQZlUl7Xou+pX0NReDriyUzN36w08yo/IunxSEtB8rTWpm
opBpNspFiaFCMnpbR6FE/D+buI5/wuyPe5oMcGjtwLfNcD7PETI2Q+UikWFG2ERBgFw7Lz1KzLGj
UrMJM26MixM5n2XuQZH0FzImCqCwm1GS/9+ZOaMwW5hQLEuIRjbVmjhm4KDPFLGv77C9yjLWnOF2
z4puoQpu1X6x98jVn/TI/VOgdx5Ihx1WxBfwkNv3dAmikqm/ui/SxAfjhlECYhdY64oMsQXZEn3L
dLzR5vay1thuBgOrJU/oOIbWPI8szeYKSpVNN5s4mp/JFaNhHd3Z/a3q6nkBKuROF0FsbgJWzLT3
7ZxvRVEd2/I4kGk4OowXewcCfzTiqpXwWwgxC5Pu7r4IC3ZojUttDbOc6+++IGAn8PV+YkiTbLaU
twZeB5kc0l7nlZ5yNTbn8TTOi1GQsb/oaafuF7xB9QV2Ll/nTyyuYM5QhcGGbEV2cit//r3a4QYE
0KwGAlfxzzPMYnzuffb8vuumkt8F2OnaOlLzsdhJTdiNaZQs4eayplzkVp99q0Wdkto16R5iTDVe
4I9afdhwYJh9MQXtuoPur+ztU2/ZkxvNzj9VpYM2CPGuGuBjh8pLyLACmFZbevhZknNE1YNSyllq
Llwya11Xa2j5Y9zPW01xAfG3uxzXQLXwjkapcS9GLmpwc6F0BAqjGeaYBs88WbDrPoCoUsUCaswK
lUYtxLPg1GgiKRS8Mp27S4an3EHjkJ6nCg9gtqMJsOmIa1DPPOwvEGYBKfnsbuOas8iZyh0K/anr
Vt3XWpfGh61CeDPZEuX60S/0Rc8bXN40BcY5KQuifgf2S83Z6tYK//j9CBvnfPiCRiVM56FO8Wjy
3dJdr0MNaBTzUdpb1FLpfbcaQAq693VWqu0szQzAmwAbR3YfpRAtKDjmyZCvynxbhQylOvmGw+9J
cJMisVYK7E0ZQleTIj/hW9E0K4jej2M+5r2G0/1jPnRHET9teN9IieX+UmOkfWu5i6r2H5IKScdr
Yb0Zb42lCBsbaddmuLCMGo4uEHtm4XkPmkRJqUBZSEeya1C9mInl4a2o9MHAbHfUFvfuFdu4pRAc
/bOzaihztLQf/+ZglG/IYgJSGTkKJMRs9iGjdblLHBgX6+/W3eupFUVvjTRlKRGlT3kbKHw5ATLt
hmKV97jfFE2tTL9U5d4q/McuX11neod+Pj+SRjwiJujET38trH4ydlevF8PsiuwoZK1GNoCM+6FI
12M0qTECbZnmVLyzh1gJKyqR7n6uB2Vsqac5HnoCPHcIaHIdJhRacKSB0MfhTku2U93TrkaR3TjX
FCYZTF96Dst5RVdobWUQ2nM9KfwABt9k8UTN3zDzGOqInzZe1KZQX2lVIoPNYBwN0/gBFWd3ItLk
7wLS0E9k9ZmlGqakAIlnwyjA5PakOlccqV+MK+xMhdQqdZcMJyMHPANsA+M902CFvyt63ba5O1eg
+ASUkkn3LCMxxwR2fyRdrfPIcP3MmLFJsfBNsovw2o2cxCYl/u4e9BQatTOheYWnSY/Ch4f4Al7G
TO9tyLFPHc1fGP11RpoOJX7cgZ0Dnqu/cOgYMa2JhYHwvJqLDl0PvCvOk4j6c3b7MptosIBboZOC
WHWqbUkJSmuUXVNMhr877da57SMWwhtyUTKWsZWbTwrdc8uJvXmamr67coOoLKPCW5zbj3dDMwbn
v62BAkiCiuQ6p14p3RN7dfBxqIRqpGRMhgtE9cWmJtEXT4hR3fwWmERnBskl7ax5BlMgSln2n7El
7pd0HHOskTrhZHoSQSbQFfGD4pxmIUw2Kshee+TISqaa48wW95kxxKEiU1ipd6dD6YAQaXNuHYcQ
KnemujKeUm4tvPFglv0xAbIsgZGtDNW8WFaSklFlLjVpYpKHBNk+WVQ3f9qh+3JEEf9Ulybsumvn
HO+jU7VlRxXmav6+mRFY+sZbZ69PnzwAIH75rLoJ/kNbJEKoIz0vuKKHyXASYU8o7yk64cQXBQms
Nf+9ZSCie1t4LfPg6x5/0hys2yB6YFnIejccEicpyOF3f0CHgEIbZy0jjM7owmUjpyv6QdwfqeV/
QlGeTbc2PB9Yhb07s9YtYlHMwQTC77EwoSt8XpUUSpqpuEGxy+eK8TykTk0QKEyUX+LBXNGlj2Z9
lmS7pz0XlqFT25WVVqZ5h4JIqgxK5UMbN2Jtqxt2YEYlNPmOWYwlIrq1cDTVGlhcLkyiXq4KEb3j
kmot/RmY4zTF0fjggUhKg2D8eE67iyICCqmq0h76vw7w4jPWJJRuqvwitDbjBCi4jfrq8UdxQaja
Gn/QsZSU4qOy7A3PkTh19k+BgWS8IYcKFT7CNWJHR/Il4HM/O8/eQLeJsbfMhcuiQm2eHmuJ8zOh
H8Qe3mnAhdTztNsYgQeBH9nEG/Kh3plP7sd3H1kStQxpDF93QS5nb6CgpLcGn7y+B/rDCNa9hzSp
sVcp7pTrQz7BqTwqnfOq0r0ZCJzbptljijmStBy9XJRGWYLAPw62OV03+676ZbVYJWWs2rjlYq9D
u66Zv5TsPesK42uWsINOeR4DyT9f0z0yeAJBgH+GZmWujTWrfBB9S2rM3hRofUXkCV4LpXjb9DQ0
WshbcOMEnFhHuCIXOHQeagGqg6HRuT9mZmkLiZjYfsUJ7h7BWDcTDVb6aEId995PtFs4QU2w5d1j
6oVmHWqcAhLnWqq11iHekVItIXD1E4lzXrIgxKjtC7bYr1Ui6k6h2EO4uiTQvlnloujiPVQBfIxJ
PO/gZRgr6EN1omBNdZ06YECTin7Yns+1SUJ849yW0tEDV4evdKVM3vtNNfhFpyM1j41qkTh1B3KK
Y0riCr6XUsOzNBjbrN6qTjDX+k+yqjBPhDq1ZqKHeTXKRmpNqPoJEVlgHpYm8//74rpJS8afzn98
n+SzXiw0Gu7aMOvyq1sQ8ZBltSpW8Stp8w+E0Op2CrC3rc2vP8hu9ZwY8zSkxiDA+r7ZtKLriDje
p/tvMPLpX8baVWk6HPCuDvUgcAiI479hdnZIpqQZQf0/VEjsh9NJ06yyM8fPBRusr8LlOJulI+tc
BRrQtFBjcP4MXAdusAUNHrAyUMm0a21GfONFTeifE/zqrS5CafXS/GyGSLNTfMDe5ZwIcCTZovRy
1eapi7dSriJgOp1ByAVkkAqbkBqcBU+NfWcIH0qes7T0+mXPcRxLn0RCU5GX3WCUi+tnzx3B4AqH
U/yaSMosUl4wPcAm/W1MdJmx9loCsqWwjIdejKoRbS40FW2eFeJkGOa9hg11lUQoW3t5gCx5ogoa
APA+TER3KdtxoirTr/2fP3vOdU2ajYxtN1ow2XNP/eE0HHmreD+q10eqElTVI/idXZXO7UgKNn90
Btl8vqujHQ9Py3gIeJBQuwqKt+gkFTiTwG93YmWi5dJCoY+jeekW9YCdWvA49/mOn5Ih6zOiJtCP
iBqunsRAf7hSIsDR1u95IJmSUoV+AzdhzJvLozUsJz4g3+kxgTEqLvuK6JBEknBD0BffuAhhuoK0
qT3mgLzKnTAK9/vGJ90GxXMxcb+U/8s5Liv7ttQaNzW4OxuaLfI0VCzbiYL+C8eSAIZ9LmE+OK+b
fzm6fPdTevAgxgUt7eGGG4WSY3Th6u9fAe6zaieANakep7uN0S8KJEIQRXzNKACOGvRoilQj3tRg
KFw9CBKyfMy0o5yC4+EkNeE8exklwAggGSqszAY1TyM3nE4875NbVaeVFXPjqpFIBzhRsK5mGwA0
5ig3wvO9V8A+3tZpDDz9t/sp5vssqrNltaQDOxSPAqXPxoHsStDelsHP7X0PQ/PsQYLtYysy+wPV
k97PJGp+TzUYrY7PAw/gZokooR70/opKiNHvJAQ3a71yIFa7BP6CNZ9E+5ndOqFq91dXos/BJ8FC
zvGYGs/cBA+azUtdddahoY9HylSii1xmVHESPzaQi5RUfh4C+QBeFm/VEJ1u7LErtCFVshLNPB0u
OpsNzeRiiRTZ+Qbkbl8vTWACsGrtUqDpEu7MOAnaMLl6BQ5DbM36lP6pq00sCpbWFUUst3rRT728
5XeL1J/TCAEI7ppn2op4oi+TFiz6MIF9qjQc5reqJGJlmNDQDp49MloXeV/0dTqpjWUC3DofB+XZ
Cjo2PA/u01iK1J/SJ5susqxF42KHS6GKM8fsP+v/2y2lWxamsk9M/DMeWwGquGnmPubv/2me7uBa
QOfeQhjrrhOjBq0XDxXSbjodK6lfC9WxRrMoRoQNU5klzCkIeVpIaFroM9IGYE8/jTbR0032LYET
YCpH3MQtAz4llYS+wTXbL7Ap0ucXaL6UoWWhleqVqqjKFE8V8Fo1j/VIe2MZEQl2PIYgjYXzt92G
Nsk7cVRwdzjJ2nGDMmWhKJxqEG31Ui7OcCSCgEKG21+zOtowe+cQQT6CAoNN6Jg6p71VH0MYmE+Z
CNaCawQB3L9VBJDTiQgT8FvpUNdKuDDR4gpNkXEX60FqnFqanWrHcSvAKrwU5mu/YIbCbkpVoMeD
sPmHfwo07yvEOmfQIQqP5pepFuSVxRvv3PinlZjsM6XwsVhjpOTi5t9752p96XxYrsIzfxkt541G
wycJGZuid5cG3dSbultif3JFc8fKP+cq9cFPF/fCK/YtbMfaL9ECk7WDcJZHTf7WfKbGMO2rWa68
Og28kephMEUKMs7Jztvc86+1WjTusdqg4JAm9oL/1eg9yAe15VMgzo1E3w9MXrzmSQN8OLYMnvz3
0TmNG+SdXbwnwHrJLtdpJsbEQtMvqnbGc9zVMKwlr+gMH72DFZsWM1IZndbV6n+bDdbXPAwG086X
vlcER8UDPlOkRofSTrT15KTNrOjMqm2SBsJg9UXXzlYcopEq0cPoT9JfdBAldCN6MzUQ8b8fJynH
eHPUYoOR5VC42EsG7GuqcYNgZ+9JSWKH0Q+DLMw9amIEIrLXF0ZWb4VdDBrRLlT3x/bwWYgWk55q
mOB62uXHTStcsy7+kFw7a/af1WPbFsc5X/UMv6laGwkodq+3hmAt1nAbt010fJYKowcwDc1cVVqA
2JZLZB3NVSaj3/FckrZADFod7GDiWZXdrUI8nzEajHCEttIUvkiHOM6FaVEta2lgLuJt+SH3rjdx
/hK2L8qzYBgxd2ypDZftC0wi1Mvuo5sUfRKS7vJIyvKAiET1QrHN2RH/24Hc56wqf/0Yz6nfN8PO
eFWQG+DepHJVn4F+1OhJH/biqmvDYjeFdRO1EQGsW/qDiwy5pnnOESmbe0x63lma9GsFuT5QpMH5
KFwpEad+2grdojXaqa8p8QYpL5qtminoa+xjPtB4JoI8zikjdKsE3eNv9Itl4wCdnPP9ysw3E5Lf
YGOJjmu5e26rZrBsdnXo/tuZgL24WwvbLXr536Y92KvXojqoxxX4kWgiGF18RaXkl4YU3jGP/9oF
ECYVW95ynGau/KChzsge39h4AdFeZLxgcKnKEOIWV3ArcBW8SYwwmS30mpNSxIszot73LsaTA2Xp
4pX++6HelHFFucIDQdSXDLxyGWa/Ppt3lqWRSUZJKraMBm8SV8VxoswifRWGsxZyixTCquK8z4/o
pWCQIK63lmyWQFwgoHpbaRFlnz3A9fsmkc/hRSLtn6kXBKLm82N/i+D65JnRcK60suL8f9SeYDPi
+040B9gI8oBGtimP7Q52/mxKdxn74fislh5YbD924rz/K0tcdI6alVsFXi69VidcBasqsreE0IXS
dgo8PMIiWD5j7OeHE7p4yJ7HN1JzoTQLeWoRUUnA2oLNBnAjRZDfuIwbKcuhiTHIQY+pJnPpjApx
z+4DcHKuZWhDBTupsq8nK7CqbD0SHPn63d6qUtl1bjXnzqj5WSHK53yrvv5lpAY+AxA+znrjjQ/x
kS2ghliiyuhNMCJbm44i9BDfap6/Ar5EKgZE8eKXrKayTUUPT/dZHrw5FHh6i5sXfhzJbB2ouxZs
NS30fhhZTCeN9Sk7qeT2Fk7jGfI4qzz+f/GUkIEfe95yBrIBIIoIb6t4I7H5vldRWgi/axHPRnoE
gTi2AnO6tbzMc6DaoUHwBuOoXsadNQdokb7lAtxh5YdPHlx+i3ftDjai4OW6RzkrWU0P7suleEFe
C9qDni2YL8ODvXsrf/BcYkV3u8m6aj3/RKYh20bUnVIi5jE18kwjIbUn7O6i8DyR9IRtIGW0gPN9
jbTVgvc0ca2RqxPHImNew8UxEziKPRdPQLhjnYE++woNNPVc1Fl+ZNXACvJmnPtCrajVnDfuEhc8
qxpmgqv3ZcjGybDB2vyiDmhPo8PSrTuyUaQFdUP3qGmhHDjC8kfww0HzhTSW+Xa14LMwWgYNVndK
kIBuKV3MUboWiU15334u26R+fZnbD5gwry25wVb4Icz7+Cgirv2JF3LmHauo9r/gM4GK255Qt2St
DrOgmTYdmpwnu3g7M5ebIFR1pbiuVT+dE7QAku09/mFSAxGUAmKLaPnIF/dD7sp+7z4JtrAiAEgL
uP9av25iqeb1C4ypVUXZZHQFMel6p/aWBiqeYnRAHQKlAa+eFkdg6kACWKKOU8hojKsvVNEpOFaD
V09bqoOdPJhK6KlyA1emKdMdJOB2uk2A5bV1XnyJP+sVrN2vvrDD1CKW/nM0vqLbrA8optuSBCsY
RHfZiW3B9uk6MfUm6tuOHqqObwjk7ePrwEz+jkedIEFEr4ECORV2WTdZMMoTDh1ufyLpHSCGLGA4
JuVcR97NOu17DYMo2Rj9aCsWEQpYpBuDiIta+fDWBx0vFdquH+WuJknCpDfDRAaX2NbUk8ev9zK0
jJrWrqaC1dYuzmdORS0D4ZeKwXoWXfOHFFw6ezDZWGa2Fyzf1nbJZ77IcMjvFXjRSUepago0PpE/
YPJGEq23JfpjzUqIHhV9JduM63jnxbLkcGn+uMQfL28IexHeUc7x+u/zNp4f34ICwaBS8Q8nskBg
fVFSsZoKFjeJmvYyOuMHaulfXjvwXpMlDH1h1s5bM6v/mwtsMyjLCbz98udtH0mMSfMcwCtaf+9K
y43wUs6VeLURqkQ2KWwOQgBXpXptZaF31KpewNiqWgUr9G+kEZNy3bOFBDbyKpUHeDsF2sEuIesF
8b0ZzwEQDEXTC7e6ocSfwoRPGgvFLblh2gcfTALc+fBYMFV7JHafQWiYk3qrGqlec7d/cGZwu0Hw
434QNWhBgTHTBp8MLLzNPsyNeqhozzQItHcFL/eDjhNzQ3PnwGNPkeubnhl2L+D/4Y2lPCaokB8d
wT4MtwDeXPS5j1eIDsGaZ5vRb11nAa2YEtOtEngzSkQRw00MUKNk+DFmVbf8zxpFRfgS3FTw9LBe
HEIFAMQMUsePJs+pXv+Mg4EqPJZqCo9kdeY+GAEDK8pUHoyOgoplq2NfslXHtciS19k40eqZdEfL
VYQ6g3u0gPfYFFV89iJQGboV74C9F3hvJnlXPfGhOD/9L/uh05vrkmJs+x14tpUHtIxcs1cfmRvj
2ClJ5OheHxJPTB43xW1LxiH2AOGGCMYT/NVKWbpDT2lBUK9FNunNYfgPPLCDtxGu0S9mM5OIcTGn
UlOWA29XgLrjHtYdgPCFv7y1j3fTILrhgyTmLC6XFCsqUR0LTPTTF35Oqrt1Btumn+GykpTd8M7t
eE4CEUgy84ICwzI3MpsyBr/im7kOQg3hLC9J5AwpSwzPmzjmB+0dqY8jcTmgIetg9nPR96ZtgeVQ
XHfKE2GMsk6KWZL2X2mDCPtPrdUVw761SFbTvw2Bs4rqsf4OUhdZYK7zeazyFbpUwprw+GAzqgYz
Xx4Rc1l5qjNJuVplgWnsWdNIwrQCdWh9BdyXJb9bys/Gr0mP3xkaKVlFfzJZ35MWdd8fawFY9UrR
FJta9J43JTHcXvW7Wxvf8m9pESsQRwljbYKQRuMOpW7kYPf9hWyZ0hXoMCahk8tYPj+U5JYfZjwx
KqLZgVD7NX4Ufg+OUx6oCsaEIvOVTeLXgICoCrxBhLpikNEBVLN+3B6GjnFuvwz79CooZ0sVlpFB
h8Xe+YT/5bYOR69LZ0S7+zMObz4zuffC0uL7aEy4rLgyDuuFqVir6zQJ9w+SCKRzi0n+Zr5eW3rg
SvGmwk9arJtLyn+vKHgw8ckh+QBRWE+Ab2EH2cpCsxI9XM6lRZBK5BSUTq5l57NHR9vtry0Rf/Kg
WrnrV+p7JCGIJm1CgFSAwKsk3HT2f+iPoU8m/+8eh9F27dDwaKbn7hFzZSlpmuuRTgOjbjBD0XeE
wYz/nrPxgBiIMtdEoe2prPzwOZPaZQy/SIbKAFDgNMpp/D7VqdocycqFz3srjBVq3XSdIEVtqkND
jbPASVKiGDzLzuCTXgq0KDKoL4/VOGj6xjvlovUlhQRTBkpuKBvEbW8Zm6YdaTk0jogF030WpQhi
E/u71qi7hoL54l6sPuw0MSyimbrQnES/r+tfBjpWG6IObbsg8pQg5pLoRbC0bwGwmh6hOTCTvs1x
EZfXqcJIdRjgQoC5d3JOIcKvVQD56lL3D+356ZK96EKeNT3rLLexFUR4ay6Lno7IZTNeu9Wi8arw
y3zXpjCfeimKNxMPAeVNnwDO/BFFIJxwCX7kuvkz1U9YWO4Id5ghwdJE4Ay2rWd+TtJST9vgV6a0
dbjDooW+T+HxH2LvHZlZwbuRloBe2BK1Sq8qV+LVl/sxwcuBvySqd8bHib02rC0ahUh+QGIExgLb
tPl/8C9os5RzlWKGEpnuQmCVYhDKBE/BZ7LXFYGOJ51gEomI/Gfyyd/opBJ5bKTg0z71SYOQ9Jua
PlndvqH4SqJfaJxGI15qTHfAHYSiOcblBuepSSYR6wEySCdKXCm4gphf73ppz0pfm3BeYEnLZ4X/
q79ZS7iIm2j6Od6NziPVUcPn3DH3y2CU77U95z99pcUw7M4iNPu6/Fv6UDRlK3w+4OHtM6yRmfSx
zzNm73rOYtlutlM8zH88uHfzaWN1h7qgu87tQAhtxF0FWrseC1CBCblADfJ0/I/d+jsH48WvNm6l
/2OwFOex3W40t3BN6UF9SvByeO+9xBkK1qQvBv6qxO67qH43QSLQ3L4ed/qfHP+t2bu9SoDFbtMy
t5tORYqe1Cmn0F3wbmhhZYSd0OoGnR+aU0sG1p/WbYP31IT9/KCTN8q+G5Aqch0TjV3UApU2Uh3W
cwE1+WzYsX3Yxv4rX64f5aXy6Itjd3y97wCld8/mjGBzShfCsD66SuZKZ9++eYwhKFkraqof+riz
Pir2FRRBIoUgiQo9P6EAv/apu9xdS8l17vvM7kR8PtO9SvSxBSaYCAyVdaJMht1O0aup4Cmgys7v
FLPIP/aX+uLBjTzqT6sgNs04Oxlm+GoydQfhgkswjT7nbBO3DG8OVmogkTLJjYFEafPnTc3bqNVy
JvIPuxVuVgLyd1Vj+H1CuhyQ2NLqS7uLj/tjHpf51JQUQNkxZYMyh+R7MrV/QFNrQoJxwGi+A72t
aK3t6rtUyNODdY88NmRsciatOCzCiQLVlcIre7nnTtHiEIQ74d9VW8OzJZioCyxrbs3BrKAGVxmR
aGv+ETg5rPs9LAVCu8IS6bJY+Bv9v3rHXoizwG1sh1b/43l+YlYB7YlkFk+NXhepWXGw9CMYpaEs
nrfaCX+j8OJ0wJ/cFd998YDAPvHq2EwMU4NXPMyIfQ6OfbZW9ZX6vuZiO9pNN9kpCjeUmKrAFlDy
zfKHjC7mLpg9+YOQuxaoxmCh9uzZ9cHNZo8XluhPiH5JlrTFo2lfiKCta8330YGGKldzB7P4laF6
VaSlYMhTQxpLgZ6JsPxfr1oFFcMwe6Zia+8xfHCR/hDOK5O2Mof+Ao7qffvPz2GQFwnwCogdRt1E
4oCP5V9QqfL4uaIxrX1oAvqy6h4VVz5GOpCjE+gMrHgffBZN2+9upJMFrWQcDofLk+UBStuXWLpV
PtavVH70NUYcf/YbNOrJBeKwnodtTZpC1wyYPIp8sk/UGd54KOyiMEZJtGV6D+MG9PUw9kQL0ON8
9G09cbX+DGIwwNa/qJW0cGhR4s7yCWd3GNDVwpcexez1rNtoD6vmgHslwsI8Brgd9TwUprBfNkuX
e+jNNR/8wGWV0flaq4YAfukj+sJsZcutVmz3ZQYmtF0exr0A8Y0ccVA/mFOOBfMXgto35/ogM/2s
Gb9aJSvpXfDjh548iWBxam9wTq4m7Bxf+jAxA+f5AOD0CNnXBoIQXIMXmv9MTLV/OX4EdxtV95+R
XOh4S7JdAWnIQouM5HEjpD4TIQNlxBGmjK0bfacQ+bA8q29y/8UAEU7/qA23QPnN9h4wMoAHtRZO
BSMJApu4PRWtjRffwh9A+/kx6ts24UaAvjLE8WbjcfWAiY+AvrUl9aJKdVTd6bdAGfkAvD7PBKAl
mhC73KOpw1wxZui1mTFHwyVED7NxKdP4z9n7mPvEXn/CYD9VkeF7MnTDsVSHCqcdjqT6miM0Hi7D
dYkrdjoZ479bCNahQVeyetEkdRWvDQ5eDev2QVnBEBkZuGaQPvAJOQNGxzYJ+XT3hTRbCpwqRa5y
eQpQ7sP2l2242VXHP9OBPqRnM02TAG4+c2sqCGZprUcwEzNdioeMpYW6frf7fqT/jTo3RD6CezKZ
3y//qiLGFdc4ro/VRiVpyjU5vfHlwM4Exbm17hU1Lk/24haA7wzdkmBiB3Ghh1h5C3gcqq+K0UXo
y42l0G3h46G+yYFs2HJvkYUdCeTTP0qvHq56EvEKS87F+AhnW4K3nwZ4oyQ19mvjghou1fJ6OXaL
esPIUCBEaJrrb9NBaSqKX7wCPt+C+mngXCCByRIRHCrI0TGn9SxQw9ABkhM6o4c+x8jGPiXu0sVz
bhMWmBumRo1A49vwCD7yjPTdWjijrAfN0gBkkUfUqeSDZsYD2oxYVdViT59vaxKzlGChfubopZGp
Mw5aSi1aiy39W95/tG20n+7u4hSvm1uubU5eWPg4iO0orpea6HvvIusonzaFdZAxyliREUYGp3nt
K3+wlpn1eXg7q1rIxHPUK4NRDhb0pqsM+UPs8sFkpruckbNfyQw+z5gk0C3V/ayc5wvz1xIj1JyR
aUGucXdkacXD8mOLF9UCc3Lg5pog1x+iNMc/D38rUZR22eH1bhuUGGiBdCz1tkmWeaAnz3Pq/MDh
iWZbooU8Xo9cCTnQ25didK8Gw+iMV06B55RV05rMH1U9KqHyTtZhXLfVn3ZCYDg9hbQJqpNi2wR6
JdFdQpBPoFvFhFOTfw2WejRfgFwRIBUOSY+ugVzbTDmt9WVuNPRThAyOvrtl9SuO03Q4hGm9aUjT
kj7Wc26EOuWrdsjB1PhhlM4C2GGFV3DBOlzlvZOnPxg7OsQM/+cpVw0Ki1yOv72Mpn9SBkJxyglB
EFfF9XalVJOyr4h3f3x2wXK/2d9tn8eF/baxfA+VI1iNYszsDavoX002msvJgcZtnMxT/d7X7LDp
T7tbW04VAtVgX4Zs3aSck0LtgvRDOYGz95ynqRcYK9xi9PfSiY5Zky8sXYN4LA2ZILmmJgvglQzy
1R93HFsWQye0kHGsTh7K2EXqfS2EYOx0quhrBsZkYffDnBWiD3OnNDM6MSs6zqNDjC+rOJNZVlbb
LlhjDA/B5Hsu60XWWUMroX5HIy8cd/jHrThqCidD2P/BbizNnCbg3CnUUQTUoJ/03uE0MEUlMYig
rnzD1Mbfin691iOD1ia7+k1vQRTLdvtl+qQrVPavEYGb+q5vsnqZBi8/OgH05wh31gO3ioOOaeRN
nVmofNESpjSyoKGMeF++kThbY4i1A86shk5ayyz22+nQC2gcfHA+IUN6+9JThpSpt6NMkZ+MTjxg
knPYrAmTgzPbtDJru9jHHOmqwTFyvmJcIFG2ndimfql8HCnupS+SNRr53gyJlw6alFyvJ8rxooqX
6NT9oH8MHwq09Vqvo2suLgv4SvXRAM3JS8xGfrslffh4Hm/idHoknwctAKr9I7ll84U1arXuriUW
jup+7og0+6ZyXiZt1MI5UdtOwTzQR9BSK5XKBdr38CjBDHpH3ZbgXSfaZiLRK/t8KR/+LTB4m3pb
APwcv+v9qL6sCFXg8fyf2pLUxpRg4gxM7SmtIndrwyrmYTeJBSW4ZtMQqx4mTNyaHVlZVIyP13aq
qmLjMiJ4x2lYHTXn23bpXKgIJquUX0xrWWUsfsj9rkH1koa+GVElSoPb0G/oeDIUNSzIsxwmPkR+
yEmJERGnueih/0/GqYFJaTUEGowCIAdYf9P4PzApomRf4YOfCaWa0EslYaRlS7AFIq8nBsHZHYnm
Kl0OtUsmvM1GOrJh5wySIar/criorrVc9ORPKN++dnh9th6IhfExPaa+PGTVpXPL4vzRVrt1s3bZ
R3nAo5CaCrcIq4nXibDdojtagZX9rP5R/1hrmsNrkcKDVZocUm2AtkDpOltWaIjcRAsuIdDZbQZG
hUOrE6N3srIgwUZz0p8EL8v7r78b9Ulgm/txIeGr4Rqi+QoT+HkzDtD1ljQL5vWBXZELGs42xTjs
qlxLhsChyW5PdbNM3N6b9nwgWtqS95Igo1pyVSkiDu9M1rzj+RIceonodtM5ISasWCcizH+nB+RX
O35PffUz8qxPAxK+11JJClZl39dq7TJhVtsHrPB79Z0fPVdOqJJ/tGIfFdOP2l3HlJfyBFCSWKKF
CTsJEn05fOm3yds7hcjFlm0VJqsXz2LTdit3hxc0z/dXrQSE1iucfLba0gWfzucYoe4RNy9USWQv
jTapEqvfTAR8WUk6Uwaw2Sdw+G7zeGX7SMDbU9BhRAET19DIOp2jzueloG8EnVftnLcZcD0MiDgC
aOsxgH7hc1eDq64ib1STIM5peeoNB3f4u7vRC5zFsK22GQU/N5b7ZGT7egvIwEHFDsVsB+LCa/e3
toy7TVFZBVbBuO3Y4OQ+9DVemYRnpGiVvc0H8gjwK3ZDHOjWlU2WbYUvSKR3Gm8e54k6XRr1aeR5
RNTh8e7dGBewVCFn4tKnVIF0eU9UsjkLSyDDynALy8gPop5daK1m9+FAxp8dRiXUzSZYiqYtSvTq
HyKqEl/pKMDpy8lXow2i3YSWR54Etl1B762+BWjtIibFF0HVUQozDOCz3A+uM3xxNynAIc6LzZZn
Bhe78ikRIEP2bPxMA8hSdIlxU9tiBGW259ASsUtAngQBlOhy3qaRX7lIH7/eDK+gQia0K+dJ86Cd
n8AR68UcNK2VRPp6li8QIDdemD4E74RqJQHnAx9ltN7cFmbcwiLGfqiAS7Fu1o5/WtDlxGiJMt+r
uz/WyxHwAilXaqMkv/o/iX9BPSV+WO2uTILmVJrLleW5x1uVNvs+J26VcurPjYPstPjzAIIMObaY
AWAdG0p8xT5gektkEAjpjBwgzdjbrRcQJha/DyJ8JRCZ4ixfcM15eu7Ltq3wgcyL6ZdGjssmoh5a
m7LQGasiUe0o5gxCVEStmhodXxJcJo9zUcmyzRvliDbbmRhQoYm+WwRH/BTzcm4IL3PPnsjUTWCB
Ug87iNVySR233+9DxfDMa7AGV3I2pxQDLwcSts17FrRznfFYNmHa9PXApZRF1ccifzw9FYROCRq8
vc1eDgluECfKJGFJqWEFdOU5fXtsfvIQGsSg8YwZj/VyK2cbeMPyeaduaMxfD8ggfW2UvOTmkwd0
Ia/2dNYK7HUS/P9vdgxgHZ/GtHko9SQ1+Ba+3ko0Zv4BOKy/UfbJB3l2GvW0p+iu4hwIuwW7HzTo
2cxFXYgtqwiKplO4Q9d+qy0GdpqvHBCfQbiJHeYy8YU/TJ2yzTMMrufTgkTGy2bdicwcvQ8ls15A
CYD34lpA6SGUx7V2j5ODNDz8qqtNRUBsGdc5CmTb6IYJs8tShP1wey1C+BvPoJR1c6gqljLte6iP
Nck3C6A635zTlHcGTgZd4fR4pd2OdqgSw3oIkF3p/LoFHSTsB6tiOboy/C1BRBBmTyI+1hcCJv9d
Exrjh373SD++JhNl9znhzzSPbHKCywC2TWMgGTVPqG9JIPxJRrd6Qmu+35MD2W5SL6uTpXiOjFkO
5V3nTN8u69q0M9vuLXYCESfNEQsi3LiY88wxbnFqMaV+RhltfZ+G+I6AMfJnbyoREG7XlsxPIyJP
Y+yKCIlD4FyyCWq31WXd87UtPsADX5JxAr7g1oC2Mp9wZ85NRUTYKFrgKiK+kMQZbXKsG6/KZSGY
1vlDAl+6aa4YPnVAfiL4rsSpRJ/kHqrKCKPkoq/kVq8QPLD0TvUyg6DDrACxhnVF8jI444xB/1A/
P8/lZ5WwkVEKPTAy/6EPbZFE1Tm4406xefXxBisWxf++BvjeKwfCgHdh8wE6O7JKgU/cgHwAwZjc
I2u3UjDvk/9TG7PkRXKE5oWNiCnQwNmt8e8+SDaTsL4/cG2DSD6v6EAu2WjgfuccvfCPe38uwsC+
ORaWUWgN563KrjHka7Z+XGcy44U9KJfGXZnW9/IwgufUyYPfALJi9QtKYfy/BodJMjW632K7I1BC
42dlaAEc7EaBY6u7BayCh5pga0Onut0aO+kCywoeYUIfusmB6gAgkkE30DSkfdzFzifnpGK88NrM
knSqB/y/r3pFVoUzmwO2p6U8Zh30GDmFYo4ujRP/T7xrEmzw9F6Kkn1p0mY+WttrK5R6LdAHHH8a
AirSh31cyXUt4a4UAaxjVVgK5L2aG4Yvy/X6FQRJvNF2EAyf0gB4Fak4HaFKcxMwJLi5Sx8+1cz6
x2z/z3vv5RGXXqU4MqOtZz6B2b1ii/MkwMlitJy++dQqK2acp5eYkydH3AtZhkWRAwJR4ywvnnPG
2Av4zLQaGpcDbnBnWtpBN510kvvOhcgUGb0vcafWzerllv5SL/7O/Gf7ebyPmQItFv46I8ynoAHy
bIJdYpfMUZhnAbbRIiu2FCNiWX++/sFvOhAVZ8KXvQMCf3v5cfVpwrgzCN89DN2cVgr+ExoBAe2i
Ahm/LBT32c3O2mxX+P7PujZL/VENVwmlS1oJR8i+zKaUrAPWJuJSclmZWXJrhzXcDT2eRJ946yRT
M/aITwKb3hSScY7MzYWoJjfmLhqzn1U4S7QxWIispQ22aa4FWL9dXmFx4Wk4DEY4SwtFANayvELu
By4s2ODX8R/AqhLmuNni3NHYVQCyZ3GDSMM5DvWm0Vk0JvXH61fYKrSfiUegXu1nmyR4u/geliH6
dMpTgeko3gYqdDk5SbAInT6XlqMoNqdM5qB1Tlg7A10crlqsmya8cx1VbeqkCaOitCjhRbxgW/Dk
zRbEcu9fnfU/LYLshBgTlMXtefdGwUfOErzH1wm60nLnhWK7ktq6YfFp0swbhdLdPVWUrmnkap2I
41FZRVdItLKGPj7txt3Lt1AoyAvXyxu+jGIhDlIep/IcIS7BNlkEXY06IuuhZb0AVnDFVM3p3dWS
GjIw8lWqkAyiHujbWnWxpCcnSjehzlPRdpxNZvSZvRyXsWf19w0R1+37oYcEFH6v47skHb7ynRJu
T3T2BHsSgU00se+QO1cpNVlyi0mFNGTs/ZuMd+lYVW3irlaHPRW/e3FccpWT53uP8PmJ1Qwjdian
KYcCg2tq6aHBEHvX602OdJSxWi86Md9u5Tu4elDknC+rgP/LxD/KX6VF9JJE2h1gYL+O0DbsGYAS
7/mnFQPVPbC8/ltb9wbKHAzT4w164KnMMVIfyipW5+Mc8RwRzQv2Ehj9SUQNEgWMBp7KF7KWU4rm
6MgglUlBbNuAw7GcfVFCTLigjIZaLxJ2M6p15rmoRYBP05k1c67P0jr1bc9hC7jxB2NERWMYBmdU
zJUDrobtXc3wGvJwXDyWqdKzU7rJtNAO6+esyF5RJ3rqvd4bMPzPCFmHOqsaHjJOrqXd6T8q7qFN
9+YMSqBZaM3vtFIdJjLXsB+WktHk4gU3dKeEALxEoOy8L+EYv+ynBj5xPSgnZwvqRVyX6UV+R+c5
1gE7nAZNpT4ah2wXJ4yGSWlEX219HymUC283xQjA1OY42ZTh3RxOEmUoKT3YPG68lRhjWiky20KZ
SuM3drWlQq0p0CMQNevmFJoWgZhic6R8iRNA16VBnH31P21VDEBGAVdmEF7Yzn1G+dYr02IjV/r/
Mkkkz4V+BaXp4ghJJ4KwMsNFItZqpcIly0Iq5hfpn93NujkCR/OosMrsc+yBN+9yfW3Bj1+CqjB+
wYAyg91f9GZUibZaN6eoaCDiVWAgwyNVZVwH8MrUe4mMU7FFaOr7c7VOOJEQ5wrwiUAivhw8zDlW
D2xdmjY6bgnfWSdBHH36k2uDsOejS9KgUdhlH8KiilBOlv+IUXwFdByG2wq+lmZ1S8TJlNIarEL6
U2yqaRNp6noMgitw6Pv6SpBxZp4S6JW4v7GKF4C7mmooHG0ZV3FLPpYtCpQ2T1axS0EbzJbyzStr
BAJxY02m2ZpkfXURm7wwhufSif9CM9tDkBrGKekX6Hp47G27I0w94bq99tIQqzx3XOYlgzlSa7xE
Zea8pHwQPixgb127g2axiGw1WoYdP0xBo0aAbQJiOO9JIZv+Wn9Irnu3t55laxVf3Br9yYy0QrEY
JobJQ/OZiJkGX2mrzXhD9KHLj6B8JWnsIsTZKiUoyL7Hu2mBE8S2FJOnXboXL07Nc2QACf7sBxUJ
uG+ffUnSqece8mNKUoyUXfCvN+nSYCa/mQMCkIzOqNXtjJEZJyPO1N+VUnNC5tgcgtQ/O06PSsO5
3ljT/fihOiBiwur29Vd4oEykHip7oVt7x73OXS8CfZ1Cwnm9e5gABRBNOC4omuCl3G3uRvGVvqot
Uox+50bjhLqQjK+XNNdmDPt2BGhI5shUlYPdlpgZMcmJ/8dpN8SZYpyzJR1LJGv9N/Yk80EuRQ3v
nB7N4DaDnueFUfVZMpGbypk99igm8OaFxdNLNJ3TAObZnbZbxBPsPiPkhtQPWTQo5VQqmUkUEYeo
pX7xGkPQJQqis/SrzZLK2ef8kIjLWoSeEJ9/Tyb9i+ZdTksBHt1hgE6emSXTo6J+x1V+4cW80DnT
+YLfX0QOTSUYaLc0UhbWRo7zgKLDYyfTiGet1HFsfjmyg3s2ggwCQMN2N4+VIZD1RPBt0EOrqDdM
opHg8zGfgiu2VEhT0Q+K4eZ8ol5fuw6iTA2AVAV35MPfsnijWyI6qQYViwgLseUkYu4EZsdvgQwx
CqAOorNK8J4pky9wLN6Z7slS4ViGM9Zz+KKuaIC8ND4R3cQKt3KTBj3xd/8ptheEXAX87g0ijuZO
BibbvLoiKSlFGJJN3QmVdMv00u4nzhQRLppsXpaG0qbIbc6b2JOf/svJ0brBOkNAJBUMrV/eMTTZ
D11BgvpG+dI10zgNIDo3jRt/autCI2FNRgvXa7gJkUBSFL5T66QRB0iKtIok6wOUXhx1gKpT5tYo
10n1TyXwSQLBf+5yTiceOUqWXVRWPukiNOdpdLlFoD4TbvnIDaThMw+0z/CcDTvfVbdvYQoqoK+B
3Q4VXypsu1AdHYvSIQl0QGH5X1QoHwmXP7pwFaG76HD0nxJJPss4OtVSMa2wcWhEcPjfS+hSSta1
dQ3mWv7km9lzYbZvsMLo8pibWkKxW4dFkQkvGdDIblUN+N6h3ISSNB59wdiboGyn+688haTYyLqM
nGIlrt76fwIEDVDdtn2ue+kzh5/pP0kqJJP8VqaaGd5XqoBvPZyiPzjUDVlbC8qMKptAp+qfdewq
v8vxD6+OiSCAgsQ4N6kYfzSVeTYF89lvJ/5r46Y1anwNhh9sCWyZJNoRfeGHCQbv5XyoYvuPlUxh
EIrzz+cAEIvmr90sz5U5GJqPZxLhT99HE95cOjEWadRzpWiNGBeXx1h8ObPbc0HWj+8a2SUFuWKS
R2gQZW7/egCItu6WxLb37Yu1KFgw3Xr6i/J0OFm9VizfJajSgTglBMikLMFl4HFkI9u0Fi/lXgQo
AGwfuTAbjCRXduD2HXltNqBOmX0Yb+fW36MHCaQ3jIRxnroSX2HEleMAowtjwSn5VTR9cpNsQtlq
SwLMgxq18++1S92cdd0FBkhRnGj+mDbjUTh5jqD8QpelBAWBya/zvbBGcQ2MDBcTC/mQNs8d2Xol
/11+G+6QsdrbrpGLgaOCA8TPKZMYeW29aTScWHE0lcXEAkGODk4jczPhqBxzLPP9x8nd0naYCcCs
IHOHgHEiUtmDC02EVLjZLu0c9YKhAWKeb6MVM67C83SLfaeaUhz2ADD/QLS2cFtwBG4H8otPbEzP
O7m9aioVDMYVzVw+ZyL8ljNr41s7kP1mcvFTGdXNG2sbqGTn+YuA8RqyIFoIBu6EtwMPkxrWw7ai
2y37Qwy+o5GIxC5m1Z8FJTY9L4q9ChfrtmcNzPQKYS2EJhdQ/Oi6c6+eaKNPumBUbXKDOLvTH8kd
hKWzTqK0mv+I4u4EUzGaueY3ckF04Ia6FYdBiSY11qnMxfvMhEpDw2ZTgjegdJD7vLk2dXkkNyd5
sw1qh+gQaAgCTHVK3YSkNkTQ6PkddUpOb8/4ADQdldbB3D4YoDLLI7k81kuoEn3TZgeHUUXeQlTu
gduIvamQvpWW+NhQU6At6FLd1qKz3AU45WWI059MvB/SyrYWVflGUjbDPG1fIYY8weUL29io0Dld
sZkGcubB0Ow9Dm8ggo7Rw7nEy/CW4pluBQsegBvrPgSDKuTZbqHwvtD1nKNNL4aq9PbQclraN5/g
CPh0QpE1ocNLmAhUGVhMECAf8TY8EKDH50LS01tsv9vi7YQN3H28spfGIa/g3ygNg+m95b9Qny0F
LLl+igr3JewhnWUQaiF9L4Wr6s1fvvooe+bhPNktbQfkJoxH+oE8VvaIiJNdUEFkv+icy8eYzscg
yEflVhwx2ye5suXtERGurg2BraTDX6ZSikIiQXNN/vfKxRauJm/V9k8FrhfNuRkcEqZzMjywxJQW
S4TGS4bFMr9chpSf9FmmxMa6nc3uzT2fEH/klAlDDzOJuM1m2lBvpua2FuzBd3wdYm2ks+D1LHei
09jblSRF8CK4moaWFWVdcg9ZLzB8Tv6s9sw3VDKUhM6AjUAkx3a9ovPY57FUBoEqbzi2LAOFKBuQ
/u1wutjSHA9dMqsDoMwSq+wEjYucpm4NfpR8uELyGQeG9om+vpDKM5FkLaU0EKuwPCYgw+B8UTjG
70UBasD0jk4PmkTmYGrfcg9RHv8UMrod0ZUSsRTKHBvwXAQ5B617QN216FLwwQRi9wUZ9RxVQMwL
fr/cGvuhYteAoMJJIvZ7UlMCxMWsB3K02Bx7OgXowRWhgjChGnafIVKEAMZdu1trbxWZOutTHJuZ
cHMsgYK/VVaU0TgjejvdPY6+I5TYe81dJETYep7agWzVCoMtkk6vRdxsxaOuu+LfwwMfLsm4DOsX
eG4gTH5Z6GJI4L2XHyXucg/xDYQr2+8n9312nIhZv2eEA/HLMwyAyIsId5vSFAq1aiJHWRB4Pb6T
HK58nztnfI/OXQ8IdtCJuKlWHB2D3tuT4tgBMQgjlzluJJf/ma85XuZd63KE81bTLPp1wCTSKLxY
e651Q6KzrrP3/s7dF2KiQvyN3qqLwFlatv5NYbW75WaMl3dUfaBnjhGXoxlM6QhDI6thpBWS2re0
cM3Ysd8YRs/dyHyFO4+l5D3sWKJ8q2Oz9diaMZcdA4WDPJYXuTCm4zDHvAVLSFePhxAJMc0D7fxd
NskWD/XPHspJBuGHzx23oNaCXrq+EGYl/rzwId95efCaC5h2DEtWyZ6cuczue8WatlKYEUl8mdPP
YpC0b8vYLXg+j5d3NIVggc92NE5WfsT/rvCfcBdswl7YxFFgzbgJtzY2Qp9FKYBFpqp1L+TndGbp
JhTN138hwzZCDmjRaQFOofofI34CUTv37xUpVGmqhDj+a4N6JhI0WzNsmWrgNavNXLw5ZFrHMZwe
UEEySV9YuSomGJUdzBufU+xbgRHnxczAlUqLFitJOrnCD/EAwyuEvRKtndllVs8Cc9ECsu7MiuA1
9BwV0uoayXR5bcR0YZMOhKkUkQN1i3y5utXN0xfuXwi45blIifrVferzHBruquQOclFILFC3nHl5
tmRiMK1vdAlQdZMhWDiAvhQ6STsUK5kDW0ONb3v7viQEONvgW/3UXiz+sobRIX+7Ys4tw3/XYIZ9
wjvw/wgTi7nQY0lQ2q6sz05nCMiS2uZ/XjXOhzZsxaeJ/pEx6q3kZp6tqMR7DlKWKCXT5oMwwdpi
uh9UjC5TAiEI0NadSIFKImrgtqPzcXFL8UG/OfWxQVTq/ic0jnXy0bhYmskhzWMsKteOIZymgJxk
NRdBNOiMU9hQ8aBRD3mfh41aXQGdHGZhPBGwlkJ8k7DXERYShBcb9TQcWD7OV0ji0YofQTMfn6Ah
VMVlLr5iWrnWNNh+4BvgT32xcN98/tQgMjdFAvKboVxMeYs2NTTPDLcwecY3hAdKER0ugc5+UO2w
PIv9EmiVZ1svbImpGPi+ILJ6k9nBXXDhRW4z+S1I+OBou5BwJtcNWQGRMaoT2ITcPDGHBK5TspKM
GbnO6WuO09TIdH/kw1mw7AWw9JxTMql6WeKKVlc1XC3wIv5i8G1tHBnyYgP6OtixF0OQ3kiIQwuK
UkwBT9V/sQxNNCy4J/BfQEj1/mTDiZktvP0o3GbsKXxUsigk7VLT/qLKqafSEVJYbMrOCYeaH7ws
f3p7e4vJW0L0V/QsysHoeJgjZ5oIXjPEqGwJGLowdb+0QGZBsYHf7d8JI1z7wucdX54GPc0aOMkg
P3IbieDrdqe0c4pQp2H9ydHu/dkriq+JuKqPPSR3n6xy0rMaDXACXr57+OV8KflvwFvzNoEqbX9o
W7sGeb8bQWiRuWJX/BwUH2BZfXUiP2aNBzeXSRWePQ0cIgIkASl4PLpXbEYfl0czOAPPSuBzPImD
wKQJP2Nkfd0hrVo+CPyB3PTroD8yXbU2bvsAp+n53H+vZScL5Rcv6k45QEIO64SFgkqOHHPuwjd0
phYR7MTUvnAk9DvHBnFnLdiy5xLgD10RxXfXEOj7lCYbuKK26PCtgaLXfJOtMi3lKgKmVst6e+5B
Cqph983ZAyaLurLImOyNBmqetd7YwCV5819G7zcfPg3TbwUQLb9D7AtSa4W+To8V/oaJ/EUBjUUk
wHWkU1p6FsFKj3qebp/cpmIGhl8LnOLuUzxHUluH8vjW/VjN3/KOVikdRbObl2ZIWxAH/D5B5trq
2nxesrNh3tE70TvjcKnk9MD388jm01tp+QykxVB6LlLl4/Eo7GA/qgrOxybW/uU5t1GWrOgVh1fA
z4mctZt/EmZkUZ53qxgLFN2lmmAIsvW2WG0M2A5si0uAOI2n74Xz68+sNF1ScN/dDi0FqLJDiAtz
a5Q39YCafHkI9wCEDwP9LO6ho9By1kjyd+N2O4u912D5NAErvHUF5R1EtPxBVqBADqH5bi59QA5v
v8uaxYh/m3ZvajAQ6v8So30Qno2xkKO2mbGY9EbUA37La79Vn8S7wjmx+mh8cajIGHVLz3UDAlzM
WBVd9dEAqkTxtXln9BUC9ctgoXXm6cxW1MgaAfrn2/kXDPncHf4NXyeT4kNJt9x4fjFF7P/rERO5
Y5kgBRV6jxx/j0ImFt3sSWe8VC397J/QrAU5I9U/SJJ/Ph3pepTiQSKA+n/HvdyA3QXGcXPdtd7q
MMTh1fM77mkN5dp2/Vqaw2pDojTrQmIwc23Mdnr8mnVVOHGU368MqT4lDGqRypKt15YcUsmYeM3K
XxlYTwZkRixn0fyi2Mo4/7hKOJkMnvJRUaBxB06jPRi1TvtLvQYlwUtS5owg13mhkyB6W97sgIER
3jRznOHrpc1y1afc3Kp/mJJikz9kMVhFmwqbdsDFxgJr2/EtOvZJ7jYhzypfOt5rFj1TIyN+8XAp
6QTnv5Ci+Cs1NetGa2QyYtjJig3vpDb73I+8Nru6FKHBT/Rt8RppUaC712u91hIvyU4l4OZngeJN
cEXyMET4gwdRpm+NnDPQU+blt/hJ9zWnGNtLtVIluRDjaPZfeQQUqEflB3uH4TB9evTTIJ7rtk4r
GqYH+Ap1mzunS0VJBLzp4v2LID8L5SKCJrspJQ8dzJfWLY1Bhbwi7SxjyQKSDaiR59g3lyduGovs
pA2tz4g0Hzt3sdxio7VK7nGJaioGkYVhZb88x5ul/v00V55rUAZi4ROJu0rNWfY8HjV1FHR7zTWo
QJ1hbI3GyRQGjMTxHSCSuo05n34ScoLbnkLnTUKqod68Zc11+ylE+lyfeaIqqi7mfe0W+yKYiRRH
53xUukjjvbJdk2XWtwyHl5ugRSA441DMqVjlVAXR9VlgZZTwfqxoyJjrTz7DKfCfzYTcrLpmtv67
nW31FnodJ9uBfqTnYQFTj2VoZy4dFiGtphNbN/0jpAuHfBILQwq6cuMpOTzwVeg+5oLNWxnw7tQN
DvnW+tcI/2gDKiRMgdNvVdz2xVb0I+/NiWt8g1Sit7eqKthoGoDhMMrM0BilnRsFJS/ZUL4PsM1E
9U3//iDCEIRnrfM2QSuavfzQZQBLNX8LHDUC7eD6MySLdk/1QyZFoHiU/HRrwah8nkVhC+zbx+ba
QWC/u5GpmY8uObdtCLEu/Bed+grqdFfDhyHlUUoS3HeWbyjYHRhwja/4MI+OpNmxdAzlVB0VNG9w
YoHfk6G5V7wCntA2hLyYKxperZy+iPdkBUT20cxiV15m2woadlM69gGY0rzhOXTFxBNlPhwGesyj
XY9F5q9SQfkhb7wKBzCrGWB9lOXQ1YHPp1asvKjsuYS+Y/a7IGe5YmvDRwrakd0PUQGXKuKvfq/c
YBmZiQDms2kJHAh70/WQwEOXPaUGsZSM9r2hCij8UecajGacnzrIyUtV5hvd6NQ8Q0cRPmbqNDXA
/R644CpBY2CUbfyqK6CUsfTPzCE/TkC0vml/42Isw3ah6FUvy4RgAskZdipzRm0C28k4GaBYKIVQ
uOz5iGHQJsMOPAf/LP/7CGrrkKFUpRInzYTL6pdHXUlHFPTUzL4t9PceBSPKy0/7gHgETcJ/oG9M
JRz0RVHdIbG3UbVFYu5umackj2uuqdhJxWl+aMOZr6XWIHoj33mFxC+2F3SVbnCbWJvUAVw5tcmd
7iZUQeFO6KqX5hfsFq9EnNq899JrpdXixJ63GvdT0dB0WJS+JeF0sIVyO4BtgmwzCxCcio+vbQLz
UuOmDUdqXIAaswhrxQma+n88mSTnR1+0EYPJHNMTSxTBbUpjkRLWX4mSS6rRt8f6uVnAOeoVoCws
sOb4dX8r5GrPgzLQr7s3UqB6Tib1JiueN0EPA+MEyfgIjA6AB9564LWd5jdE+QOzPFzIGhC7poAv
VZbC4Zxc6nMv7jcPR5aohgDDdn/RWou7mvN5Hy71OI01ZpbgyER06CKQC6+RhMKaIA3G93khY6DP
A3Km3PtBst4ss5jV8Xz66JXEiibqGtwDf1DE8u7Mxm7AWGhe8zLs1sueqqOP8ybje6DKrOzQ1q8J
ENWAKyLz3rFevp/RfKgitt6ToQSBXTVKfIyspm9uPJlhZMGAgNepE7FP2NHfkaydp3wRAVFJ6TAT
JfVekfAv6Sa7mtUK+KWzU+dtZGdn3OtQhnTi/sM/VA1oEz+x2btFWh7m4uS4Jgr1TPcfHHDbR4EW
C/ibgO1MQD8NaqupIJmjwhkURnfPi3hrwXDsqeu+k9oy9DemzkO+KIjAMcbkFg34GE9CMCF4kw26
BhOOc4LzmHvaQCch4rf059Fjvv33FkYRWkSFhGAMhNrQlTBAKWQdmee7/uDk9vVgmQsp7oqvYu3z
GE4LDAMMlo1S9OfEHN6mjGx0kYCcAwHxpAWhgHH4/dlHW2KAwpf39ErNRxaEbdZUXTShHPTzWgXV
mGCk6cbhqU1gPYvYasASWp5rysYXe7pvHwvAyOeoGpHL8fIVBGgWGmFz6kpNrOFLMUx6R7/iRxqu
nhlENOuZIFG3j0gk+B3FlGhhntzffL8FVUZRnSGVY5und+dDjos7Qmx7WMpussLvw3EAqdgsD7ty
CYen8JoVPcLAhe3pP0WBwwcu5L8lgoiyVOvIphcclkGzQ7S/F0Vg0a3IcFDvn/yyIwI2+AAjQB3X
GSW4teJ5olKS8C2d5r5wEnCyZ5WuPX/6q78Y+lgMHDY8mAShfAlETCRV/MUAorXnUjuMNtMNZzW8
x2U8m70t6exDBhGzkal57fiQMwCwG6pSDqaA9qHuSRgVZt3WxHhqYwHECuf0kvA8mKg998Ay1c1R
4+C0Blu60Lgy8xHh3YwSnNe5539vaZ61Ca1heF/R66liU6E6FRIhOI+UI/sV3Ax2IxfgTxy/a955
/JUyhJN7JlCUXEBXRev7aeExeiMYNpy5u0UXz7BW4k23rf/a/tameiScJ4ODbUzcxNKi7kL3hMs5
6NTBEjErYS8waJL/uALyyvA014mgVAwJNOhLEGzkcMB0Cs9GNQwirIhCP2Pe1imMRm7X3lLxmw9w
7LLAIq3j6ZTBW3pybzEyh7ui+/daCB1SFOGuO4K9ajVJ3JlFdA9ePcZDmwX9soeCcX0pdO6CBAHy
tJzm3iclre0kR53/OtTCgOdWfN215MmQWbFgH2E3F0Q0Z8PvfYJXEEc3tj2apBOy56c/31Qz4n2s
XcOs35X4UBx7C9Xb428jf7OLEbkd+L77yHnEOZgfpK+9zyja8hZPK4h9J7/j/U+3VhX1o7uXBRcA
eaMKTuO5T0XXbd3pkdPd6/0KUDioxXVs/g/db9oZvsIQXoaaQKCP5ZXBYwn9zAxXdWPVNItHu9ZL
Fe241OwhVNVfuoas8yw1mmSRj9UjZ6n5ZuJgYh0m2TbFjLDERxD/cNvSkNffAfnhScZL1XgyGgJR
Ag/qLECEVoj9TXIAx8drzMK90bET2oJdR0jdldxuo1tT9o2r6gbbCzUzW3cArAQkdlv1EylzgQgT
I407MsnPTQwZZlxXV8Bj7kIjnh1gaH2hp+NoRjxUA0ggL8Sk2ilABdlFaGZbB8U0EAQR8/96S1cC
q9mkF9rYhT3Zv241YUEdqLorOb2YbD8IZsTvOuBBfoeULU4850N9eW5fOytrI5MuyPWfKWCSWHG3
DDov9vGGncgNraEf8ff9fKlat5xt3nGDyKp97kURoRccbYjd4wlgYT7uovXvWM1+bbS6n5SMsG05
9qGkT0mafhkg4UFs1GVq9tNouw1ucRlAgM9c2R6ALw5Tj+XDtoKtIB/01PupM7F12p2xa43Y0Eg6
Al2UOCM9rY+g1cVl5STOouSfsR5NYzb+NRYr5xplS0D6qPpINbLjxLDk2Yv2lGdk2r+irXg3YJm/
nWRh/bx3NZ81gOLloar1Bd3GefPkeA5sThY0Y51kof4F3LZ+brS9NDuWBU11eAHA/oiyDmUkG261
Kh45kBwrIc8xv8ApP0rP+DbPRSjbTE7MYRn3XE0+teMitRsaOyfB2gaJ/cjDFHuQPvIz+nSfeh/i
ZHeSLaOSHhaNwp5Q/10nDf/GN3BFVwRGA5BuaS0VGlTxZBPJHESYYJWKQRgtSsVzc6fy/m82gnJ3
hG7fq3omfGhG4ZCbOKUYgZEcQ3v3JnaucrGFnLCPV6CtPVNrCPmtwxxobDhDiZoVGCywZmBcykY7
yEeDaOjEtbt95HgPjlSLNNy4frvDlD1dMYI1bS0649E/NveoC+sW+m57teq4ScOsOodFuuVnc3io
BfIW0vUJ8KC+WfX0AADJgSYOLkFUUuBzpXAsICO+9VaLzFcj8vjT2DwwmrzBRWhiCqRcW5S4R9ue
ortt1I1GO0au9wf7YzDTSLFqz1f1Sa3C+JqUsaZwefl1rX1x1NVhTgGWTawWekG1YGBau/db+2aa
nrtlvTmlpvL/YvYT1FvEy84+oDrJ9xdkcRlj4lIjs0+ACRUZTarzkeVH4cCvyonBkLas5nNB1+oV
3tDH5YfAHuxVbWt8ps26NtjyoWskqE9dWgRNAHSilAqqM9jbJLR+E+bKdimS+8w/I2dq9JUCA3qv
yEeXFjjoSY6xM3Y1Qb7/8wHYvx2ospqw7Nj00gmAnVYWKX4l4hoYugySv+91t6xKCcFcX5Ote+vo
m1+BXr2qA5/NAFNQWsE2M2cJpihlp/iujmHBy2qFLCWeT64WWc4z0rE80U4Ryhjee/FTyEateer4
BIpEVGTzsnCeifDY8e5lrLPXoQVHoFuzS94+LVgUEiEYalt6eetLY6sVXPq9cfZr9+/oTNfyGl6X
vHiOIM/yH7E7Lvr2bPCwP+jSHe4Ld4CnzGfBMcRhGWeF6yap2vm2Ztj1E0yH4wY270Y2Z5/izUxm
GE/WE8G0+Z8G2iLZMifeuxH9j7gquFPhQTKXbdrSZhpcwJv22l0Y+2kJNCFVlIIvqNi4/Qa7aEo6
JCi5AM2JCRzljxTP1k0e68HlP7cRxG/Wh+KF5O+lNXpAZdKw86+Pr89pA1ZqzpApk04x/fp2TP+6
BCRA7gwGo9n3FXzh24o3+LVZOcFKvkqUPmnMlSHN/E3GZeiO4vfFlD/5iAN14Vr6pjjoBiC7FqZ3
YdbllMy6X0GjjHmDsD1gN8KH5CN8nRSqrYa1yRBnJYf6jGCtH7K0aNfjgG+Y3tUZYeLxpg66cM+v
USsrU1Owt1FnK8vBpUHr98BOTHUpk3lDu80aHeWmIotmVSAig2uOt6+lU14DTgrOVq+cda6UoPlF
Eqy2/akrkKeaMPfLYK42m96xo/wpj0lQYDoyrulO7SMY05Wn6C5TV5jwMYDr8b30irqTF2NFzX1y
m9gWhR0NyrWBCaIbRDaSIhnHi1wANP8lcHn90IqnFRFptEFdVxTauebPDLM4BC2m/1WTzn65Y41O
/aVN4FOYglibXUG0roRK7MNDZAs6B5U47cu8uVDY78MPfOAaN+sJ6O1H6q0lZRiM/q0zpOejcOmO
SleqGuIh8RjzXQGbSpnRSc+Gng2c3UZvbBQRww54P2mZpy8cArbGB9iV2CwTFhXPsZOVWrvgxoIH
EIaNXYePi1okEvkrICkaUGZTokS3WeBxAsA9ZG6G3ge3CpsyQ3FZ0LL3KuPG2GDL+dEZlIzJde2R
qIcL6Qzi8XtauA68ikFhBNCIPENKbXAgloL0D7o7D2jbIiIZNZxqS5bq9Qpbap52GfEOuHi0DLIs
I5JDURLKLyZLJl5gA0fT1fs8eVQP/2mL90nHF/YS/M+CZifCJ5TAemUyUb/GeNaFUTFX6Zazxlyz
RC/GHiXRQIyLtCpf34hlQbGRf8SHEM5Nj79YMKAps/fbOO0ysITcN7o9dYrDUog/QYIQWq+SQHPK
LXcLzxVaDUydxW8ydTVkw/NxUJ0lcdPuKkrph1wdeGDdz/mox2bEH8Q6bBVWiZjMLA2UkZiEv8lU
kuq+pmhWEHmFwIDigkF6XMchosNpu2iRqyBbhTrqzHqA7tdkiBD2eDc1eq0j7NN0BiOjVNWXgoHC
tcJIsBM/rsBHY6mKVT04wCdXPdX+zpYj3dKlk0pZt8BzlXwrf9oIo8ZR/YEA2H+yeGQkVjY+Oqv1
BdbOmM+BK3yQmq+70MBbcJyfg4vLq5cUh3zTTjZROTKOqvw/bcA8+++5g6iC2uepMrLGniB+amkw
onwonGZ/fRtsH+xjFFU3fGHdAZXaFOHHb3RAT4Xb5wTIyRIJ2fQAo1+U+wvfApQoLYp7mOcXhtks
uE/A9QRx6NjX3rD90AwQScPFkaRDJ2uoZsN2lgEI8AEaa0ZFgnmtEQJ8LpRTcLCN9/QoQLI53W6O
qs+JLb01heZx58O0nI/eECHVEcmKarv+PUdRq3EItL+1Pjnn8UiPu9ZzBe3VjdDYfR+a6i9qTbvL
c8xdQ/ChuSrs21w5pNg/5FlL4Li08Llj0wV8dDK81uT17KkP+pK2FG8IQe7CBTPnbar/2KTfkll1
SOIZiS55jq+nLa08g68l6ZvLwu9Idip826gyLShC5I04rH5nv3HZ7l2lpI9iSSYNSO/kkLIJ/fnU
0LqJIeuXIgT57m2wnHxyYfzU+TuVXcZDHwySdqKSGmonIY7NDmFXNIilygt4VQPOWR3tOVPnss3N
MtU3PrA9Kje6nFBnhgLnZxM8gJknovO1GEo7FSfgIOVT6yg8nD5Gg079NIZVHGOvxyXSHYiy2CUq
0d1fHxvJB0e2kw6yUKvoT1nydRJwqWjq/kiDbcgtACRSIfd4Q0xaORyfroTrLxDNnwrbq4lysGUd
ApyLFNWLp70GyeZOZGq/u1UBuqmAFbdwmqBtKOwqy5eZYVBTuJrSHODfW3cJETkliKZEh82tiUXy
380zussScjziVviAPbVCvoWMq90dUlv7DgqtYoQbsbUlhnkLMG8G7jym0SC5p2wezVYihiJG3jZ7
OT2fJVQ0P4sAJM5Eyz2o2reysvtFjTiBqz46fDCSIAMVYp9iDrgsIfgI++60LywD+Unp+ZMGY1Os
O5Pyo+KI3hmA+nVEaf4+E8bxIRGKUdBcGvVVL/gSpAJ8/QZ+DafiwuvzZL6ow4a2eOSdrUjgjjDc
3q6O6Od/Y6cujHDA+KsA11A+/giITWwUSlXwav7TRuObB5+nK/I7r7dpjRf0hnK7MwuAglwOLeeb
ZabvZKEqqSPbFXEI91R9X8QbKhIQCJHSXDX6fiAnCj667N/sD3msGOnQ97jdv+Q8rvUuMicEM0gC
ch20Q1i6VT9AareuK6QlxNd4JKEsHA8CNqIV1GW6PCFTwkcXZTm2ebSPRreOpOH0RPfIUAlyiDzT
Lv5stl6ikJLTQ3qk9MJmLZ18jb+yV3sq6joBTegdClVA9tUolqS2KkYUEEXSUENIOa9XAzF0Z+bM
Su5V4N41eeWaWKscNl+AxG5VqrfNxItltTYM0hti3h3t5IGY2c+6RjIBEPhoMrSuh7EDAhgXSVqY
jGqxuwpi4rwD7Dj/CwVZIV2UZ+n5bMgRIN+SZI+WwWzoigdhVEb85oNicjNsvNXDZNcEq5UIjrhw
Q/fBTZ1wOL40YNCUU/ujpu7efkDJfI848PB9YpZ37g41FaWfXDKGpOQZFBT8bSqlKVH9X+94HcpN
FVnwPgXEk6LuHZt++ucLr3Pdy5dZi4dRvDEzk4wKU1oHrsNBaPqce0ePyw4r6ZKLsYCqsVPsmNzh
/cC9HSfmIQePXwJclyJbgap4qdsdStZbNne4fDAVr5RNmrCRceN1a+hyq4WyD33aGJYp2QUwNCl+
dEpapCAGC2U3xmXlXs1kMBMyZZzH2Gfmz8wmY0pEY3ZFfTthQCrfFzs7pyWxfHyEEClnR4TKP1yc
z+4N72scI8yMg+9tO0fXjt6CpGsXIeu2E67RQmVc32zz+ipiA2kvABpASNs2tQH79umAp0pF8cp9
/htECgtFONgZ8qjYaQwKNYH5SXiHLmFNUVZgRyFbgFRkM2bPDEHuGc54eTnchffW8wzKjhPk/i5r
p0LLWWSrwZARO3Tauj8kzYdvR6774jj2je9BFrhb4eDTGwWbySfYfjSg1Gyr4J2fMm9wHbzwgj25
V4Il7Wfrl9/5/oFOnSEbWYzEWqKiYswUlwXmcDAxz98OZNFacZaPah31DKma2p8VDpUVoWV+PiyC
3hVKWZcpKDZgm6QVgrpu6PVUoxXPZjgXF5E7zrVYvAd1xppWFMPFzT45/Zg1NlOkYFkjLedW+cDI
NEZ/SeselVoG7blggyLkTLapeOmxg44D0imquPkD/EUHay2eV2dcMn5X5HT9MHfyeIH5kMT1oGkV
D2jLVviz2qhP3Ry6GcBMomXttQNLe1Gfgc8wRRMJGXx0HmaEmUcnbR//xRuXHhB4801me3h/Spar
7Qf7T5z5zxGaBuvpe6JVmpMboN/cAvr957NMqpuJoeKmh//RMOI6ZBOBYaggluvmG9LjRwBfTyIf
5kXH9IQqy8yXquvZ6SUfMt9q/dOmCBBKm0DVWrPllVW+aKIjqClzCuHmmnLpzXGGgQ57d/QxRJQQ
33yocti8W5jKJ6+QybYxgI6SW6vsIAgGeHjcW/b1dkCFf2eTWuRE3PjmULj+LuOf95R5PWpDeKcv
fEfm5xFAbWByXAl0n8lLecBlDKojPv0WBkJXNSp2pa763TMcWgTuybujK3KKq4HEBnF4nkPhEa7z
yRDy/wso7lLPXnkHCEVGA0D6KWK1vlOTzNtw7SIjObTMlKSc/YQZAlwKBwYyAJX8KPDRg8G0qp3E
CgHLjCtZNYPRpo7NfwjS9DllyKdfsSGw0fAmRpcLPpZgIgqNkUJPKxhxuyfEQB23FQ0MGjP73J2K
EgnQQkL5YaI5FLR/lhwIW1kknMB90UX4b+U50oO+XFh41H0toynl/PMrVOWNRQV56ua9YAT+KNBr
lLUc1Fl9EUOf404RK1X6+LoTEAAFejLgI+oPBChYOMj6LULBLq5FU3k6TTbi7Uu5A8qeCOLYXUSz
OiLf3VlbJMQB1OOfK8Ok6usT9rnXWhmsXMD0XUz23B6pixH0qnGoM6TCZcSChUkaFPvvp3yKscjD
TKzz119gYrdfMGkHNairjRZ05sqRpXkCFaP84Ki8GtXCpMM71R+onZob7b0KaCaA2zpR7pZx1sHq
jtihINkNgrgxQtpAurCl9023O542Ps7OsZSN5XV6VgYN/dnirdapUMh3nmDoSC8H02GZoPBEH7fC
UWVpAH5BI1epTiPCyyosfrZlYJuneo9fpkO8+5G8Ays2XizvGx3wKv5MAbcyeC4QCaLlxnbV9xjf
pXGoHBNmCDL0oLawiGe9deH8Xi2y82fUpUobBOMljzVbkr8PqbbdMrQJ6ZVsEvBepRo3iSNT8pOd
u0Fyv/mB3mH32FBPMd4iyM3xzOPF/hoNgRyRYtuLy9Q3VT+i75fIqIVsfd9hLU34a8Cc8NxWH8ay
QpKKhlOox+aa5pZt9FotQtemkUsNEMyFFk8//iIMs5IkwoLiin7oF06pnymEqmYxSk9QVlYUJpYm
BbeDdViGNffzYYXbzigzk2cfIDmtnMnzTWkrue4/iRk4myB/ejfKWJKDIV7IF23p/NifzNAj7tSi
oMaqruNyZHBGy4Dv4AyXTKqGYcOnLfTMOubx/NMLyltZKi8JC4Y6DZha9GkuLzVtw3G5OJTi5m4R
fk4FFjZjjFw/Sk0xex7WU7RIan96qStAKttmUXuJaD7uqOcoxy5zZe85xRFJEJ8hIq0fQFqloC1o
EjLmhMxwIPG/jL2olIZqlXVtwJI0S+UAqwzESYoNJdTZWID4tQGwwDxNQkmjHQr2W8R419UpuCO0
PhX1IQQvxOKBayjvl8rYUk12Vpm0txxQRHLFtUKwDActkoMpjBfUvS97oWyOFueCk4uf8X/iYC7Q
MSIf/lKPuOsZYBJ5J9NOco4UMoNZsY+mFltcrhfzFkm4vcP5f8vFU2MBoR3sWt2l055YJn4/7F3h
88uh0ohjC1alhs7ifnU2mKLe5VlYOw1t0dgI06cX1iS7xb6+xZifw6hKokE9eMMIFgMYSa1c/1EN
PXjuiBPtS/OGP5/sGwgPJN9MP0r6Q05Qow9PF3Xbnt/Sb+nYeI+umM0UxCYOwVt4Kc8utOYx4a+L
x4wHKQM2zhXYEunZhvQkYbbbhPR4JgeOdUPnnNTQFqxq/HDfgAlpHuSsKPyp2W/SqOQl1rFAC68E
LcvNlvbPEK+2DGwT8+ZlDtDgHsfnuHO1gCWGwoGdSBsE2V12qAQKXtK6FbaNxkJtIbXd+7CjYvK/
3Xmd1nYoLR9BXKhCFuzWP4drzG34VzF2TaISOcXISdjWMJ0Hao7R6AVvHnAw7vxQM2G2xLiIPUil
bwSQE9PtwBQn8Ba39uSYGN3B75li8G+CQaVzjFAb39jGK46URfIpDwwUoft1p7kEMjQQduFg8TVJ
NZHrb+t75H0VGNHKLt1Di2IjwBDkGciCiBDONqxeWNMiVOwDcsKsY/rOgnxjPteQ7TRMa4uEOEkJ
aWn4NNHxxxQm5kpmnq6qQfFK6Qds77ik6g45f2R+YR3MOtqF/4uJcRSCIzyo/uxsASr1hX6agTt3
zbsKweiLMyryF+m8wnxlbBpTPpXyYLLkra1z9o0iNGESeTz85EokX2k+ldmDcYTiB5pRQktiAL9w
UORtCttltYne03DN5w6hKiYGOXVbQHoCSas5PcA1+L+phR4Ua/J8ieEH1j1D/hDlckwMJWGcWBh+
wb9STyN0nguJExygUvScpS+W4HFEfWFzva/QBco/BNob8egQqZ6KSv9cb0/pV0bxyKq75e3se3cE
Xicln3ZKK6SxuYxIQqkWbVdXm5iJMmzpg5WvEvMxun5K8X7DjSQGkOTcwQSXxYIatD5qgVZ4mDwP
XmeZlO4PEsXPXn4izvV8LyQGkD25KR4EI24QIn3SXMeLuFE9JIZ1DOLhBZoI0UtZfVWJDXOgohFL
C66BpllAYla4PEIpA0C3HyIDC4AWN3Os07AQhpk+zSzwI/Ue88NfdLuH7o/G12BqTMe2sm6kF9ma
uw/c7AYlszIUSr9OEoOFgX3EBUR5RLX0L638W3FvS46B4IWLZmC12qnViA5CxcHmPiFw5qv9ms+1
2Q+l+mlEiuVuLY3juLFUee1vFoWzal/gGz5VaNjnYR9ZoikqdrzNCGj2uixv2LEMqJ7epFOrV+I3
IBxKW1A7b+3k19AR3ulDZXcpzP+l8NBK3dUHaW6OMr79sLQ8evaI0Is2DczbMvT7UDkhKLoap5u8
bj7XoIl1LZAI4GOe0CKRS1Y9XHeQUXXoF43Ok9aYiaKr0yIvaQOL/blO+VAcqQQ6R7GETvgKCG9H
t3DmbmIkXQIqIxZQT2MsXJWgUrdbWHBQGQKjSGvquXnsZN0CLIZUYb6P+Q7y7Gy/USluU3TNj6KH
4Cld60CE+0ZP4HDWNc0Agx5E2rHKdqhB9RoAn+2Yj1AbVEzi4ErxUlNqM6GBF4lp6qgzn7hFPRbL
Dr+btB8gOCpLitYrRixlOgBpOkcKGw8dhzr2UxE1C7nIfi2ZBoDEY2FVZ8VI/MKw4/IpX6pNytSd
Jra6Bs1XbDdpzcZW/oXVS7225GxlDiyAywOXXCBbmG/AL2M0Fs8yTd24DPHev/5pICfBSjrFgSyB
NSiCrICrC0CID5L4rgWswcGMu25KQIxjVUGSgBSng/44hBGyb1yoGuAp9zDuN+ntR68eFgE105X5
8Cz8xPmXcc38GLin427dzU8sCSBiHkH+gD2Ty7Qxg4HV/RGhwP0lZe/upPzFttA+skrQjMSSngJy
Ghj8SXMNRvmI8mHpUT0nbti7nZuGEpTxrflCeo4oZPncs/aGZ0vwqFq3OoKxq4a9jhx0Makq8CNN
LN3bxbv/sg2dkqqQ/jorYU7HdMJKbZi7+o3Qp0MBWzpBCu6d1unqD9EkuN8UgWwQmbYqHCsUerUM
aMthqUyeFUYlq56EZiN5MKWpVgLHRq3YfF+bDsRfBbEcxnEgb6URbnmIk55Xe0b5H5G4OTcuiQCY
d+8YebDhJjx8KwjIm204+1r62Xt/J8lSnH7Ms1P4cC9gn1phrqigfmG/UdHDyMUvTI5ayccH+YDE
7QnyoD82Z2v8i+dRGlV21cI5tUJyA0hukdn5DHWvzJ/vp55XW1gPG6oubtcvoSTACJErS3H2Y3fX
E6vKZOV81Fi3woKoQgzZBDaUsquzN4Z2UXylA8Tn3C4SaoW/1i7GvI3gpaAVF5BTQ2FH9ef9SkgT
8YohagMLYsCrMhU8bhwDtVESasdoI4CZpa9FJlUY04QSxp/BPTFB5l+r9O9L0h79OewEnh7uR+5H
j4hakwYKw6ZW+MSXuJFBzy3fbCBYpp03z4Vn2W5b1WO62rKxkOPs9HH20Q7mWVFjaSFhgMtTGaQi
qkViNth+aiq5PG/gfU/CwlRH7UprXh3Lx4cvaEcV4/XJced6ub+znjHcwvfwaMNS986pblWcBnQz
/3Y5vZVQqCUzSk7ul+qJMxXfXwTBcvSphpHuBInFLLcSjG5Lp+VNqJLp5IBWUG45XB4NuA1t6EpO
8n7h7L5D/A8bUGko9mSQZH6x5N7BxcygoImYTiGydVRk1pe4Vx3q7v0VQfl5VLdgezv7rzOL5U/w
Mbxe4/AlUpeXHmJOZif2ZbKp7FN7taRNT3GSPjfuvmln/HNk6RiUxPZNVLpt7ab55lZ8fRtqq4PQ
jHaBYSdikVJb5yd6hIchOAjCe3I9dodBv0ECz7+1S3KOfzvJJSPnecbGdPyy75eCO1WQlr8ckxGT
tVJ1jr5OCC5ZvtURfdTchHWXC/qaujvHhrAgsar5KWgUHO3GZjc5EGT+xqj3SoGTc4YTkg7JNT7L
fSySy+UbrQ1/ViQExrlZwXCU4bQOc7QOW/NLUHSZoAtdC/FSNWJc2kh/mLmb+pjCCaRCjh5i4Avz
CZlExsA123ly4BXtis8vPbU0ZfOP6hy+PYbqyRJQBuAywng69vWQbXY765KUl131YIe5AKDmTvaf
TVUtkr6PdK5xb5hrWiB+SHiMR8s/LVxMG1sBjwRKDJZKSaADKLXJCFj8zykNEiYLPjGIRTo8Wfft
wo8u4yI9Nwgt7ZgsFac0hwW0rE38bUwZl6OnZ6oLBhmIGsmNyCykbsgAXjntpWbF7y9tdjdV+Px3
7obA7ZWtCZSaXzUFUiX/a5E8A8NtHPlg8IIepRzALQEY/VIRY942or5YZn7ADx2oBjVPJ35ZNSLS
G8frPU+/JyrM3nyrH0gRj/ULaAL103jMip6NbGQteBStuBu72qaw2T4UhT1XpnSZhvMowaftnc2o
hl58xT+LRqcnMoarmJg487IMGmCPzIaRPt9SqlfJsqkWZi1/Gv3qVDoEDfBL25JurZDPs6BWWxE1
Nv/jiCwmL5dx7twoiphNFnmMzNEROLFXsVulxPhOGG8VDzh5pitMkGnqyDf9dPjH4QBVAuvFMpb/
pnSliHXMkUX+StVrua47XT+IofuzUh86n5zLjgF3sjLiyc4vJHEKzhjqE6sXIemzPDw7bDjwe4sR
uUqAx2ws8LtBW3ndExfWeYAOAzVHhSEE6wa5g7Qo1Xwxn2Az8G3Mrl0yM2ao32P/mYbF3/OgF0Zo
vAva8C+MK5sXQQ3iu2hRKJFqfWQnh7ucarepAZzB4z5yxVV8yiSKNJQexYZhCYeHD2fCXntxyAmD
31JpZHHeIgiCilZUrGohaUJRxU04aipKa/oZgn7phSk6KZWGkcn1jR6P0iF8bwyBsE2uWnjNYqIU
WuP/a6zx2fAJiLfoTygZjcKomGuzyobi7ywNIGXA5R19tjeu9B0W64apW9Ow08Z/odrzLVeGaiC9
9xvlxozbDWOHh1Ki6d6bcqTOe5nUCSmKgHckFGfb0q7eOqtChIvnxANlRfMcEJPb7CXLq/0SXogP
59QULAoCADvWpqO+mRMWKaCtXfNAAv3jid1c5nD2AEM6n1G3B3mfCt0miY4pdfR0VSh5dgHrxJ6h
+PmxX3tUOZDrm384iA8xYke1Xoy9tdhbQenVSLhyPTCmxJEEKsgiZAmom+EX7Rt/D4xE/uJnyqih
KofOZBF41YqSVZU+YXE+Er3dnDBLr1OfndXR7Op7Htw/MKwMosNgf4UF3CYEuUEeXDi/dF7hgWrb
jcSMMlzhNYxLVRs1ooqTuJFV96a5L1XYWnE2a3nykVx18a60GmjI+KHIIghi13brOnSTuv7sn3oT
7K4J6kDitevgNrLvzrfr3JYqp5RfC9aKZzwTkybo3YJlgpU7QfUFxbXJZaHxEVQwXPsrLR+wksfQ
BlbbgNFBspS2GFl1hEpEuZ6+JWyQ9QXnTHV1XmzAPPaIlW94AwXILD+jUnf3bjQ1Ml5GGeCpp7HZ
wGTLX6DkgocrzYtdDBSf8EotSXKMW8mLXaFlJyg/dFOCREmGPFrUi6rPb18DOu6Ri5P0M6wJuiP5
gfAk4Y7R4kp8Ii5xzlvVJNYYOUivlRAiUfKSoCYsJsBynRucsCpp1+VhF50s8RPOlWVRaoexU4nL
sChD2XiD3GeFCa4poJMACxV0SKwy3slvsKp6cBiEn12hSW1/Fjl6KTPQywMSp+hbNV+P5HdljifC
Sg5MmnKI5BVYPWao85U5Bjaa/nroxohi0IsMDbAkKzFsBAW5x7tmaFGazqgptAQ1+9V5h/6CVhXC
EgkyYXRH7o96ajF3gIGYPEY5OVxIUrhEwOZrNZ0upvyVyqKhNg+e07FSinqqxVqKzPiAYmRbqDyB
WZUAfJzy0Dnqvrkkske+pQzZBdsffEmdIHcUwfFoxNqiEUZ0LLHkuTQzpkUC/EeyvACti9Zhs88d
AxN2n98LzqTWJp1UeLe/IGoHBXI6ZTJWaYO0yfxKdpEIZIsll370aDYxSwRvLCQT77Cw+6bCeRCI
PnEaisKY2I8+d4pJnnc/bFY6cpfy8JP7n9KC4O/IF0O/zHA7AQEVhGHVROTBODC+Na/cVDp4kK/r
fxBkBUVJIN5x4US7tix9nmAkl0MGWRj/qcyRHJonmNgFwUAntIKAWiqTpSYuFrMJ/AKMrRO2kp15
9mO3MrYbPgdKHCItLEyDMqMUPVJtqWmVRO3zXmEKgFOApNozwbRbqbSFhGgMJRThakxa3pUWLbgF
u1Nork5J75jxRoLLjFJutXVWa1TuFfpRG7puHloj0YT2fZ0fBX36V6Mt+cqHttJ5SJWHpYqevedt
bWJ2GwZdec4t8bw5HSXWuq6SknRqiyEyMgtt2BLX1isdfrVcl1fIyZ71J2eHHTt+S8oGWgjCVM5R
qY4hABWlwV/i1dRopZMd9nH3PCpQ90g+o3PepItSiWAQabPQX6GImoHO9yZ4vdwogseQUpWiBubt
aKXbTsdPNag4sH0RVakLD/OjkqMRZdAKeanFUwakoH4W+cJEdsvEbNGeFyFnDV/xNvUiktDyXQBt
9Emnen/+S6/KpKtQHXF0TAvqrZmYilQzJS73OUDqkj5ZXuvCj7hNc+Mu/fih1WJ0N+l7P9Guhu73
OoAOubnczyU07n6zBt+okfPsEnuprkBk+KtR5r2Mbt+SDK8tjXxSJKNlVj/K4FkEoyNKgu770XQR
yTM7k6i1h+kb9KcY/fuey4b5kaSxSjTCAxzFMoe55doAOvNXDt3ZZCkrsl1TkSrLoFvf0Y386rzU
hlPY01aQFufiab9LoCofj7/gyfm2XIBOteg6M6fcUuFUQAArHvWquBH4FQtxDghtScjEBm7djj6u
Fio2sPyrloCSrMucnuaWL1zF9vH9eDORvYFJx8qkUKeZThleouDqo1kEnZRjurUKZwR56izjqmq+
ykhCqj6FEY+1reptPpVYJeMLHGY0a/iwJAAkvxi73kNEapdY/KaOKEd9gxdWvCBg6zNmHMZ32c2M
V6FNCnERUvFGYIPURG1jlZP0I4iUnSf3Z8Ax70zTIMy/n5zXqbHD68p31geVoUYVku2WDvaI10On
Syg9/Kx6hJrOuhEIMG/7FosSRMmmJIEUbAu/wi+qYCUF9vd+2twPkuXdQJx4wSoR0cvyi42ebEJj
Q8q9do7mPk1qiOQ9SIqVeZ4fwiaPE5WqWVn8aWRsP3yMMgCpDRZDUUWyZznLEyQXefEOTJvwP2VU
veQqeujEvTSN22vJhw9wfDeggBP3JUwdyfzpihACvJeEsBlNj0qvWJpgJTQmnwJlmq9WBAoYJmfP
jwhBjeHswoEztRqDGRLJwYHPAkfpu1wJs625Sn/G/E9k91pbvwgS/6wMA/9gTjA4OF3N2FSsMU51
NkoJy5TjR7veu6rEK+aJ+rnCrx3wXSmZtfGFCCwD9oiLUaQB9un2qg2J3oVT41xoT3z7BAnKFmrS
gekyCLAORjn5XqrSUaV8bYYrMkpcldAHQLDNkdtRGKGe7ZJZzlpVx8JzXHE+A3YAoHtedOF7XPn7
Ok38ZuOAHcI4GsMWImqYHr0SYfgnklEYOCWVuHG6fbYArVXtQVInbso/J1GeVpXpCeWFzDBIEQPw
hzmsf/lBjpRVCO6ryyHwvZclHy7spE0NNZ9G8CCvR1sqHzXMQD+EaU0AKC2bbwztaqj/xklyIMJS
wtKrM3ibXAuJQN4dLdPOaRICfAqUat8fAu2/zMb/4FjObxKjjqdq4rYd2VGjOTknyqso+cMsRny1
LG6y6buoWzaZwNvxgjt9jPJo8B37K2j4tUloHILgQwXCWFwwATr6fm8UIOHQiLD5Gf+8RjZVmYsC
fPXFB0t7eNCJ69xXSgkFZVEop3RgLoW46G1/lpqekzmAtkIiJoJhg0O8JY3VQnNYuhbIMkH1bh5w
G/D4er1ORG8RZu5jC1HXplhJaoYHdoi55cHXSDo2AiZsAp64SmAY1LgOF8gUOp1nTyqgcUDFUpO2
PW9BwGanzSrCvgsrMRjWpYaAIvR7QOxCjnqXo+iAacEcbNTHMXFwgGf5vpGbicMTXekz+4yzReZt
5ezy+rddx8vxjB7qTp7smKsXzbjpJaQwJZ2KpcPEF55OtJINcDJTrJg5PIRua3RCpqvEpjRMx/e9
eXRL33hCmBTN+YuUzyBaAaauavMNZ2N6W9Zoj5aTQ9+SCPBodqj6efQeG7ne1ELuDLUC1Pi0Z1v8
PMsV6pa4SQKNRL1HLWTQ+0rPso+EWPXdmS5W6zFp9SO5OnpJ58NSv/SynoQ1BwATm+0X0GXzBoel
zT/Jj+6uY1iSIFoIrpgn541++u3GC0YO+V9O5zejAqkG+O5UtPEahbiKuYe3o817KEM2VbEaON+B
JZ/FmAWXTKC8HK1eZeNkZ6sDVe75ZWzr7jdPz/U1xQa/gWETZORsKYZdBnORVud80W4ZmhCJ3dyS
mrmM9b/wNDkk4Jsd9gBdjpdqDs0J8j0sO0fDuCcN8o7RxHnOBN74viSDfA/kSxmPVDlGYOgtyK3w
o4GYKPCcztp88bnevvdSobb3pSibJsoA/nQex/98bxyjtCapSykPWd6hXYSK3T8PDzK/AxhcFtzz
SeOzSS4xmIuAbwBtMAgbQVFBIBXQWk7znNkR+Egs2JVY6iYm9F/yMLGmAwn22fJ0iXQCNGHfKHGm
oIy89kO/HTR5eptPsnqLdQDblheGZK6fMZWfkTPKWw+iSH1i1E5z5YIsWuJ6PqBXTkIfbbvNqA22
ud8mov2Pka06leGwAa6wCP4NQrXLjmjznyMbW4v5wfID+xZsuijVY4+nw9zu5qxY9BKNUqGjYwex
CanC3iDmHU6N5/AARFvlj92cg3dpe+qHRBp4363PSfzACtO0XiCk15Pkrq8564BmS8YfSE/nkcoX
mlXIEr6HMCh9XWlw6QOj4GCajnsCYE+NERqqIvuCSzwSKhxwq49eyAyUI7ezF9hcYS4U51vElxJj
6EXEBOJgQAQLkCWcW3qpTjMb/4FmOBzXjxSuk2f3FMpu6B0FV8xusb+xHf//qlnFj4PQY4LYFppZ
hI1KcFe0HcVKF6eNR5GsfpsxZl6unBvydyuJV4UDeZCJCmX/fJxogoB/q1wa7kDmHokRow51hPFs
ZD6J4YmxRMrXDbl1aO0QtXCmpXfMNvQVtOl1sIJH8wkoQKjT+vyEAwl+86wsEEsrBg5KyDm63yXa
qjllbiFSkQlrAU+vqLP3DPvYHd8oX8bnY3DJdzKPl1I3qHFtmFzxWttfj06ReGzjn7h87+JYY0GB
EfKPYIUJLZpN7g8VU6RA02q4gsP8MC/bs45m2j3rFozLQZDvdlo7dp/oNDGNgWSHXOP4Gta5S/8u
XKBOFlbqqLvTwevlQ5jnWxy/0MSIs1Ay684SF6vL9F9ryDfloXEM0z1GGl/zBPcQQmz0waeJ//Vk
VODOh8+WjrClrYV9prdDd41dYW5KBHyiG8oDY1qSIVYEP1TgvmUQGFGTaCHwUw2+FF0CBEU3tkw0
7PCqlEFzCk45xIs5+RG81Di31O1zxTLWMnqClFtvVbCyQIzs8Cxd1PGtls0AqZTTcQ75WC6oiKPs
CUkos7QifaI9rGhVgTWA2T4pGnJgQRXR4qfoQeJ3aJ8yJNsN9VsoHmuNbTPHBAOxwCspwoJXtc2B
5punp8erOytUJWgHGeVKVp9SNxPhxSz0IxO7OUSIwOE0ElnfTcxdBpCojVGfjoe6jfp5oAoqZiIC
wQ39Q4fTZJWucpv9mmuJA1kYs31TkKKxFdMoMQyj8rXxH59OzpbBMEoteyL8C7QDhSUOKfayBguv
FMRJKHIrzIex+jEmly3GY1o9+d3gQaZxAhPb4JSKl0rbuLy1hy6O2oWlu5xpepnZ8KAZFcnL+pci
RmY3NZZ6CaHxkdha9U9PJjsGoVT4vK9T1/hnc0M/DMsqU2gfp2l0Ub63w1bca+ReCvBLoXfqPBk6
kDoXsEsSSxTggfLhLcFem5Ams3TufK1J4Q7GDMffL5WW5mK33Mu4raIoDlpNSeIdEaE+pdFnHXCR
V4M4wIiYXt8SJCUS0aVpZNYHLUi/CyTeD7uE21EegO2acUNa7AhEDsxHy+ACLvM8oJGepXO5RI9v
sFXHJYJYVnpBrbhHFkVXbTsCiUe2nwzSSjgeNlR8008zjKPzOPvHOjkO8mphyKuut8F8lPGjlBUQ
LM5l71c9BWiNjl9jkYEbLQHJNu7Q52BwdqZOQiPJlkuPeqV0WLWg6Zluprq/BloLh0uEUjGWkamt
y2uidCcQtnGIwwfbSwJHx4GvY65iatlkQCjYOaWPtdz9S/wJWa+9eVaZCNvun8RhDqQRWp/n9Fbb
1z1qx35ZXqwiUpu7X1xzlp5X53QgT5Z0V7AQlN+rGGKuCoedyjfyX4LNb1krFkvRdL4uI/F/Mfp2
8HoYAzen7pN7u36ZenuLntHcmWoRxph9GEeoqLA3TRremqqH9y/GbgAlDYvy5p9W1+0tCn/DUg5Z
qc6bhI03NrAFkiixhgQfWJ0fUoVPCkVSDrM3o9g0KDkhClMx79VJEWF3KQKxDaKHijT7xm6R7l3v
XLsfhjOBOWvKhN1TKSZDtETS7Ngl6Le1uzqFW/41AtIk5UzV1xWpsiNbReTuT9spEyv+nUUJQIx9
TvcLmGWGbdeL7Ymxy28Sk1A/bdvPC6YR++14eUMw1y9moXyyEY7/Vlwukbjcvxmg+1eTjDXUmLWx
OKP3nzQ8d4ZJ0Loo8Rxx+d51GaotC+sdmF2rUEUu7bE0wmDhrHdlQao6DO+dmn4zklElblNjx9ZR
iQPjjNS+wUy1xLUfNkDFl360EaBLZhG4Ox1QnxY/fb3StIPZVv8S72NXlhdwvTJoulv9h957f3vN
gy5qyClj2OtvGgweMbVWlC0GAfByvQzqiFS6Qmu7oc5COQU0LQs8Iu6aTAI3mW/5YYYxOHlbT94h
IP8S57QpGajp92XwD9DU7oVOaeKX9O+VMlQwdXVfgO4eIk/ROPBkPlntqZWDFuKOXNQfz/9TNb54
nATkaxiQ8Pm670oCeGj9Q0gNyV8volRRslX9SDOu32AbPtVAvELdm0ydR001AhBO6G/evuGGI6dD
ZiQyqg8Qh+NOaiX46sc+3GIWdvzZ8a80qGdmk9cB/gYjRVHWnpPOfg04o/Wv5MiXCUdD4051AOjI
gLRcKs24VSl7i1DD9MpRiFVVXjSVzpelAhav6qzIm/1e+YEGw+dv6+Vo9EM4W3nkCYSlHEbZ7at+
pdVaDf7EGvUU+unhI+9dFnnrvc+HJk6dgl4rG6pc6yh8RzWIqQu3Mf7ZVrbdwCyb9cE87WTxYs3I
H48feN3PooppmKtzoVhV0YMEPhWTUZXnBEdhTIEye956wMsM6V9kpUelPx5vU6PTCTxv7VKOxMqp
ovGvvwjuyuoCkki1E48RmH70QnwWSHNuQujs/DuDdgakLnVJi2d0oN4mYzyVOj1pHkIa6s+rUi2p
68jRHsyf9Jq34o4mWuh9HuxwuDxXmRVG9TZwaUNl+sN2hoUBE5ytZcKQM8zMxdanrlL5qXAVLyJ9
iIKOSYKtsST5k0pzd+kO3RB07QiyoTmOsitompKAS5rgdAn4UGKXWlyG+MFhewwLAHD7v8hzi5T8
fjWVoipLZnOLepuzXhBBAHTjBwZR5SljDZ73Kr2xdJtz4rxvjjlzcehywoqVWD67BSR4R3GSDzEb
UhMjVc8oWLEbxCN53VMIJq17blddDg6HBZg9IifgPq8VUxyoPJiMqqtUo2ZeEMjCf7BBO8G4a06r
Xx6WS7SktgwDLuMJaPJyv0JfNMI4LwTZ8HZlOYwIYsQiO8ogBsNF7QzpMdAHIdF3dXPiVF1/OYkM
Y0UrXBIpJcRuj/64PrY/HcdSEPulwZ75BjWz8nbTXB4TaBvxCijegdYy2yYAZiz8D1pQtVbkqfV+
GmYIWEnzxyZqFoZvOW4pCkAzX+bJuIuOpWfAfPH7KLUAMJUiKRRFV70joeR9SPUFKa3vFQJKpIkK
efvDVsA38/z3ic08TIXDKhVvgvt1BU7HY0gLtj93t4paoEdE31MDjT0wCkEu8Qam5D/b99rMS6pF
oxvGy+L8btJX6TYhNqMzCfZDV0ivoUawN5/yL/jVzcX394VKztcRPKHmTvPOfcgR+Zeh7leus+K5
y59tuH3ddOgpB4D2WxDcHTLQPtKAuz/jj2cPHPKs2d2sa33aY2GlNJxr0DwDbBGhJ0xwk3DpUuia
wJhXaHFcdHTCnY2GlP/SVurPjky0EcleCZtSpBubIsPNyOy5vfUlP+XGnKc7DYSvohEEApQEeRIN
yOvWneRp9V+c8mvuyKo/uGkMQlrNPC7Q4WX3AxFlf2vPWxZYqrhH3aR16lQECWnqgGHJrWye9bYi
jEFi9o31nwDVWXNMtS4uEAFIuV4S6Q3UHcBnbdyMHyuCiKaxs9jqTc6Fp9/MAYbvBKbZd45CYvKw
U1qQFRYzXL40Lswughwpk76Bk1zxRIolbFWx+Z2euzGjX9TUNYXncsZLl7XZZjqA64v3Sd8Bf63r
VaJcWqksmkiIVXqHjA/JW9MypvbF5fcqS4G+CvF00uk0HUtQfmhcUL07r8adJZPhfulnMXKForW6
dWfJU13c7WrM+mqoQvPWZXwWDNUh1RM/WnfTEpNGEnayic9fReLfdYHK3rjZjMwcFvT7zqm/GoIk
WDrubwr+dPq1KRklVQmTvwNZ4sxDT1C6ZnOmNXF/IJ4qOAR7nm/FHukkY0L9u+j2s6/nTPG6n4Me
qKmt2CS/a2p3MvM/GWK0yL6VyyUXu2M+TWAeMSm12VwGpIzzP/jD7Rn1DV7kiI1MCdKP+OdZqYD2
RKkcgpe727MERbBYO90CRGFI0gOV7a2j0IsRIIofxkshi7knDWz5Ib5lEKalj6uBKyqREv4DIGEq
1ck4EP4O2dmtUYuAUqO/bDc8APomx1LuZCecHNH5YqcYvpeWvGzqV87mcbC0O7MkxA04r7Z4fkvl
0dAvVgLpNgptBem6M5q7KYnTGKn4aE+1sNHJt5spw+eINw++8juYE8J5quwYGVwTSUytcdIICD7a
5BKiDO3a5UYrh0fqY4LZKvkB0Lq6TomQe98+04WDopsVIvNI/ONLiWX9NBDJABo/9pEKA2UEN3E6
2Pd5bUTO2jhruabE+sbkz+VDKxeAFKpR4bu+mjtTdl0NbjdDwfCvdQFCEpE8dLiBN1w2yFwJGCEF
fM9VWwgbhQqGuZ33FFpx14UbYyCap0xCm+NM9+LhRIcxS0pgZW3tzrxJt2zvKcjzRIR6izCMYVVn
MkP7dBnG888U7C1+dg8Zh+z2NsLN2+cUPwVRf1tKMFEjrzugwOK8MpZUgga7o0rNhbeSyqlY7WDc
TyAEgzyebimwg9uchzkQGehSM8h8mh/Nmn5ugG/5OYn2M3tiPkEeLBWukCvzFYP8elRCzKUdxM8V
0CwDL8MFM7lR10aCW/urcOx9N//xd24oXLlwPdoVbpWWrBT8AJmKhaHBeEPjVxqMKKZejgz8mMt3
Zl9Gz4CvdqNgn8DCKehkwEBxPQazLSqGSbNlS6IgHF443fOXAmnXCZCXaj0qoeCsDC8Z5FU+phId
uWaIurpGR7MP9kYZV6O6kTE0ggv9H87Tp9x95acoH9rGxZ0iaT1Jb1asgCbKsOZWVayd0GDKRBPS
StrpwK0HfvZvySBHwa339ffE/vbt4obaLm69PvL5SaLJW9DDIYmoX/Yr0j9wnec2WWTxErIlXWhq
NtBGYS3oSA3QaYci2EdxxybrpCHzDdg81fbG1H6yy68PCnGD42k/4AcDpEY3QWRYY4lycm0JsZQl
PqKl8b3ez2ltNmtvJgrwdj8B4nLy90pXH7yaMw1laXNOB/Qn1blQYIIE6zAyFM3r5+iBVrAGHMLG
ONcRnMhrI+jU8utLgYztghiWBTFRzggdspG6ANcdS5mcX4oVUaoxccfOSsCOm3+n2EA2OSOX3Dgr
xoDmvvLrluYi6dy/rBtgE0Qs6G/syBpttJSxLbj0J0BQcU1pWtzxO/o0drXAYugMl0V51RSkZcXZ
gs47Q3l1GZaD6DrydMDeldO7VERTRWesKidsCX/6taQGz/AtSO1ZS9rilYgs375B5CuIIRWDWY8F
Dlh+x/ffzDeR/ezFabkURWB9mxXkZqNE5R3mvoR16dLAs4tOWBfNTgTnoypo0dppTupFzcmcRiZt
vrSpKyc/pIIqaxpSxwyqzzkySMacGmTvZcSHYnrCWXCBrKO7Zs//xf/56qSYq+9cPYaJ9McXjTUb
dWmdj6xkhirPednKyhWPHIk6u/gcLfXDBLrvQ9XIsJXQbIPvLW3BNBioLzTVaVHyx+tm9A6Ikj74
TiHdL8GICOH95xHCeCf4kBOlgjuSD+iAUDuWPr08mUiYnOVaWuSnDI/xvIUZ4FlcYejgGPKCwoTf
pXHPrA7i1ksxGSqtbXei+HJzXeushHtgRApTm7f82qFhotYOXe+4X5xPzWFoWesjJ+frYp19SMEb
Qs3VFUqIvymWcPwlYpEu5eLvu+VlD93OETy0pIhPgcTTY8KF0laLkMYROTrieUK0eUH+jDgib5DM
s4DsecOPKm91wZ835ewmr2KPtLlJ6qAVSul3HtwyW+iZvTvas7QK+riybsLMSz2evauFlMaaRPsM
82tezOeoMIKDi6busQp17f34dF5HsDCKf1XCILgenu2CmQzyLbulkhhv4zXPj7wDOzQG3vgiYMS0
eMnPTJLpS4roZKzuMOnM6hxY8PXEc4ebiB8YBedaSqLZzQ5TO9M8+Ca93ou2y3gN0PnFnADg70eW
OzIRoqagJlv9pn2+WLn9ST0JrYAKMCNUBTgaL5G+7ydtwPJoHLO13ai5t/juE2ktksxMoiL/FdSi
Wyf2/QJ8VLEOG4/uCCpvh4QdcZGjI7UasVgBf1oYM0pSrM+PsfxXb5tYVqXsim8dEH3owWyFtzrp
u79JaBTgCaf20pwBLx+F9qeT32VV5pHjKfzCksUOuoc6hlJUGxV7CfrewmZBmZR12mtovuovSDBH
ogrYD5xeKfn1Zn7FJ2X4hduFqJmGCc1ANurm+TidSvvg3wdbV1AuUt7Z7RFu9IBHwdVysekZqCRI
LCWV/qgm/9OT+2QVMvKwfx/a5O/XUHWabgQL55Pp0oaaowonHZSnIuN2jK5+VeMxPtXvBjXLwSPp
ZyneJ4J70nxip1P3ALqNNS04iTMPwUBbVXaTqXCK0H2FW5cOrj351jEUUApbb2vxzRmRRIjTj9MA
dkgMrAzDra7PTPlEeyBAEPP8NtMMlq2C72GpkrTPxZKdK+x10P29WaRhkpn956MoCTrbigFJ+ldo
5Fn3FIVJDoNy95lKGFkn3C76ZIhx6kmtE46ZhJAQuhRXS2UQihae6knYCYv1UVX7ruYtxBnQXVud
wlsCebq31YDafJ6EEL75dYNZf55tFGJSDRJk9sl0/+teloNgKSQdykChzOSTZKw/gPnVn0NHkIyz
uyHiT39F2Twea4JGSvRpnCAfw1zoIuKdOSQKKLDxCU7/T/AMAKGVHdS0dnYaakX6FREWT2fyL3dH
Mv2aZm0LIUeiH/7BtsOW1QTWf1dF0ughMVdTIJHk2ONaIKUtVBdmJ5Tg48hONIc/ZUQ/dvR5G8+p
jXxybiKOz63KyPNH/QwKG9nEqNFDYOPvkDiTx+NGKcX8PAjV64kee/H7b1klftglWsrOVPrF613l
01BJOH8f5BcywQEGJPFKy4ZnmHy0SFwNHjZOhzWdus0kyQ9zVbzhdV017AQtv31pVjryukyAGQSF
cO1V5wmKB0iY+N01JF7doo6Cwztk/qbnlhRiAGmFD/uyC/NTbetcuVIJCV2su2uXak9TP6zrxAyV
VibWB7dUQiHqC9oa3prY9H+cdGpy/Dm8DZFBNjqGKVH+Aszur+APjWYGsHBF9QJX6R40O2jPA4up
qRQz4PdvRl1ucdTqGc04FcDLP82TDqIUZ+K2q+/UyfhSRLfqvm9PfunDXF6d/8nDCn6q2TMWlfRe
NKBKG/1P1xWgrvvJqxWkp1xPu+jt4YhuIhlkstvE/kpbAA5sxF7eyQFQhIQqIlnT7oA2sAnN9KFq
wQpPiVq7do/gv2OsSgYsFyy6bF2fGCV1aTNrPnoD2fjuN5MkSGJFeG39Ym3RbVcwvSD5sfva4yAN
S7ui7NWrC7ePU8pyGIHFcmFbTNVHhK2rw3N33qCyJclRePA1V0nMAJgiQF2BCrmhvr7OHqlwcTQI
JBUyuQSkuiSzzSLWhUNdt3h1AEYumt1CvxaPmUZUNrCII3CQM+PSiyTq9C9TnzARlT48W945a5Lu
gOST0NxpGtbhQDUzHeOTOnJ2VklOsf1RZugPE3d9vzQLsoNtUqLQdHAY8flRO69LJMa+LLZ0yzMA
4/RyUG6EwKpPKlvamSm1hEyS8rXaWnPetGx0xA2KGzv1HBww8APSQZgkS11g3gJCB3jOMSh+jB7I
xPEGEa/4R+PvW22Ss1/M069NokJLPYn3+5/Rle/ELnVg50MmQyPge25yDjUoCCEzMoVRD73x0kZW
ChVzIkXFC7cT/CzsmruSSGGdAqCsYUHP5+EEA1k7rWEj7Sq7efzNFI4geVuXWSevgQHYt/BmYdtM
1VdcGs2SN1CaYh3216Q/DT4CULgI+ZtTsTp73XRPMdneYIwqWyoJsup37h+Z7SmwInWWW1SKRYE/
uehhr524Pm6IriPor9h2rj8U425MNwL5QGz1aQ+fwWlX3KNYTYzvZ18q5T2rTcI14PaVTHoXA4iL
3xaKvXwAYP84im38NGN70j9imoj4+qn0lDSsL3/y3VeR11aKYb0AkpVw5Nn4q3U0lAaalMQFTDtM
IYU68OYOQvy6st5DtiaMNCp65d1CvBbwRj/SXTcWyuEtYGOUF2liSGHjYFp4oLBetgRCMmDmRDHt
E1LNVV1crl10HgaKuuDVe2+jrkc4bCCpMgVQwhkraB1S27irHJgShjx+unYOVs0UtQPwfIlRRtv3
fD91w2GVIfp2oYiuf5E5HR5EzaFkZ1/pN2T52dwv3L0z9ZPXNoxPuUMGPI8XNCn3CRBRruSn/AFl
qM1W+kWWjKDboyldO51OfDlgXE/v2MKZod4tSUfPvwj/GpfkMPkPy9CMksTHxKq/x7rc+cdG5dAL
7ZZFl8XMeZq90cqTi+NMbnpuqdDHC6A6FZr8/bpAM7rTADO7wW8qVbDYc+4v10x/UCYI2jTB+Fh+
UGghjtZwrrCeizp6NIWZ4WE8npdMKXHaH/eGyVD8mXWoO5mN3XHnvO8WoI5bQkSHyyyNCngWJoPO
/zDgynmsG7qPxamdsUsKj9ig09/gqlXNyx328h50UDJdeifnvyozn440rPtm1bL4Qn94BAzHYNR4
UrG605SqoZdfy/gy4JpT4KuFi9F7EWS8ooZil8epNeAFkYtj4c4wzlZzKEWt0usJIODMxiltOU4G
Y+oLxhqvshTmaeyOImUTEfUJD7hvxXdf/2QYzIlcmdI3U4yaUKu/OixzCaQew7njrpqCsKgmZzg4
aEVdk0ONEsMqp4+GcT9gd16kml6i/PDn8Ca/3XSwzbU0qze7hGB+BTcAtP3mSZyfnpKbDtRRW0kG
itpCrImUpZfir5vXQWK/EhLRCqzX7lguxl9LYU9Z81lQF22/rnYnoOD0YKYpNR7G5j4KHNX1HjIG
VM8zQYtPTFZys+FBgrJXqzAWMG6xq7yYdVyQMZ+kcOBDiX+FdSziVKhwrJkaaIDdFmXkZDftoiwK
ixb0hog0HkL5CyOi3n2ABJqrFoG3B2OfR+lXHM/nFyxJzrSEbIFTPddmFYsZQljvy5ZMLa4u9kbo
ShamBLXEeCh6qc1G4YN2PWLsGxAsVC3w6XQ7X7d45nOoOVsfpioJ/kqIOf0tlNRruRyvrnxHIYHH
jHJhl9j7hcPi+kNJ+PDbeUcD9bzW/OavTVrB9m9EzegGymMaqyzI6jiFy5G1ru0OzAVoh22vMtIp
1HV2qzuskgGuxpZUwEo3mvQqLJplAMJplXIPEoTOTW399hHwanOjjjze7+KNk2iffkhH4QeWI0/C
SI5VTvpCw6zh97kGlGl0d9OTNHLRsFyIL8QlSmgZi1TvBrKqttPRJIZEpBVeReOJQhMhRN/PfpTn
8A477LEuZxd6rFCJXVSr0Et4ORzCQsSqOLbG+IRQyoq3w+61R5oLZQsW2Fki4Zq/n6EmcVb4JI92
Deb6DPalZDR72i1ZKcENe3TWKmVc1/qstn8l562GBp86mfpRaJVhU0jCC2/0Rmsk1Na7LZRtuAqF
ZTsDi3ga5FwRbNca+dCccdBz5MAVYgT4eb5KAe9UTWabnAI0CFx3/iqSFoSSnR4/5F9uAW59AF2x
uSkZGXdJugGARchY3DlEH0c8f3FDjN8ErN3vD67gZRriJH8L/6wlkbZael1ETWo3DVTpLww5iueI
TaXXzORnHKqtnPmpoVMSVxzdQnHScunHbDtUXhnq3YRMbd/JBYEV63AqAJC5sKTUQ4nS05R+oof6
zM1gTpApHGOtNHykp0VmzLKBppOZz+MF/dS9QzLxLxHCMQdaznroDO8vJ78fb3xF5ml3DPPN8V7K
/8aN4RYv2qdhdr/GJApnefmzfUDiqzJJlBW3/+58HSgqlo5Npc0bgsY4rvDXkFRkfo4elO0H9qLL
vHzf/1JruvyoqAxB1LPBc6M7AsdD1g1q7IQ1eZKtPb9xpQjbVISGHE1ftxEcavPqLcfpwi8q3XKd
xLaa7vmUD1syapsETtlqBvvq9T40FPhiT8V+X27C3ZkZDRBe5jn8byAFcGX9SrdcnuO21TFYJZR1
CaQQ5+Q+7dtMr7UEVwTX6OvGebADCCC1NA4HPESId0W/MyZPQ7C4g/onSY+KKdyGYU6YUNowv1c1
9qlWO9ku7ZpJahH09d/xVSRDsxhRtruBX+9QW8BRotyiRKsxTtdTDy/Nx7oR20fLkbXq0SVIzHFi
BOr1YynkTgoFUiK13gtmOr6ZpVp3/4AKQI/h7HziFHcxvFLTHTE+Qj8U7uT33dDuF/0rDXsOJ3OC
VmoNtshVrMWfIAPLXzkQYEP7/lsCEt+4ai774pGsOyD7a75f9D9Dj0URw/IhsYY95gUgbmT04QMX
+rJKrY76y6tHUmRLs974P7vbt3d9w07cnoSDYIKv2T61oTY726avA2Uh5RwrqFVh5tXeU3apr4Ok
NOmuWq19n1Aldpp925p6ROdfyKR1F72F3OlRPd0vW0NRl/enaP18mC3rYgAfmj0LXU+RYVAn3qoA
Vz+j4GtriM77db/icLXC75WTgLC1eU7S7bS1axSOj/SH03YwJYV8AzTO+yYkAjwXjQ5sUeYKinUj
7ioHubsHiEBTYJIjys4dVpxov8qjQvkUTI9xHL4dMghJe8dmqxZsdeaG4siunPQi/zEwhrb7pqUn
f9wNO60bWMSuMTdWT3GgNhs2JaOTMutDm+b4WbhBMtmSy7HNUdf4hosdAEc6YkPw6JfnyTQqycB1
lz1q2RjihfYwEHA/cJAGw0T7nLNukOQ+riI4zkRrHqsg5ybaKQL1cnAEVY6VDGAAdGONojzrMx0w
Qysdu0S+RY5xM/C3SI9gPIApNTa9rCnW3RTQgne9UvX5KENicAGIkTJVK4zk4gDankHiZnxbBBin
smb+yMWvwpAgXnfSnPyN2gA06jhXDitxwXhdGxb3At8VjFu39fSR87qvivh5YjqtXOEsSmmYJIf5
4H9lQPoa9vIHzsSr2CULkmGGYEL1Mh5J3EjwZMFanLsyvKwtX1iFfDoecyfLeAuXMVdI3efOx6VP
40XCLhJaIwejCvfkAZrZgMjBH0k9F9cAuTGjFje27RO6kVu/TSUKWGlsby/PCj3c4wpVfwmYLqFm
yXsId3a6aGPD3zrucfFe2S6l58hsxtl3FxlmW572O58OwsRPTlMBNbDU1/DWKRTejK1V3QrEgrwh
B2pctscbfHXnkLgmpCG7gEKyG0+fheRdF3x5p11DxosRqV2j5bYgv/Yyop/lszI0N7dGB/d0Iy+Q
GY5ZfspGdRETlQw+M0HP+C9U4XfHPUgGo5DTzDoPildUO7BVtsnfL/GP5bEQAqZRU46KJcOVXssA
U/Mm4ufAPxprLjxWj7/zOPyNrs0PtloWGCp1k6PAS9niYG61Uay1WcVKaRBCzul0a8u95ptxwFe/
KWTMbt8iMoqtumcl5iSMB2ceADm6oipM5yTp7rSvy/j6elWMTGR6+MxwE67Ph20qLKxlgECh7Aei
J/7LsmGsZO6wuOwsbp1enz9xNpj8tv26KHtVNghFhEUUp3tYaWCzPR16KWCgW1oNyhnT2tcF1nSa
hfVtmFDrWelDOzWspAMn7D3TyvqebDxFxn01svBJYmOBvxhOmIL1lYjMye5Bg/9E/1GyYewNVLt1
o7KBpbOCjMXz9RWJBqVAbm9xykcpA9AqOPQ5ZjQRXQvjP32VwlTgsdSb7aqhPFW0vgXHqCmJ+WTe
TM7p0Dy9t2Nea++GeVONxwInQQ0i7yrBzTYVil9jRr9SjzQ19cxVqY7SwIwNMwNwGDB6lTUJ3eHj
ELjhadqXjzWIuAyzNohAXtyBadmpAI1wuPRpclyxz5j9sP9Ieh28xJBBRkxg9P6gc7CdpPOuzGM8
AOioU02kG0DXMGdiz0/Qx8/Df/ht+RP4yjMAo6/utiPc1ijCG2K+TuLgBEU4f4PaBztvde+xf9dJ
5+Y3WmvUYXZKMe1WfB9gDzWgQlk9ORXFa1JNMKYSZX1XvPCoJV8l3lb9WuWOc3uz//6G2dQrSdGy
wbRsP0ei+phZLiVL2o4ErMItdGOY8ISaqnxkFSkzN6xzjBfVpNtrBcB3zrdxPIoOqq0c24SLv1Bk
6SHhJdIv6GiCb44AhlZ0BJhuBx8pOz+CKiGtbQgpsswK8iI8JRIDyy/FuLvczzGCuK3ogEN4/H+/
4Zcbu4imlXq4jiRuwsXCnfzgccPy/rWpXqax9519VHovde75Fq35df76/ozBVXXs5aPpj4Pxu1Jt
Th6SyaPjDmeHOLVZn/9KW4vHZ2dwW3VryvlCbm7T2GUxzkBVW0oygV7CYl8JqKeNPUZ6BahBgrSO
Be2nvqdwjWlKrpoYUw+MKM7NZCLX/miBPl0Txpkmn48rFrGvPy2JzcP195FBni3CWP0rr7Z66VAf
vs5itmWIUBhr+8JJ4rXMn9fZhk6wL7nyOLcs7qyrMw5uOCosiHFCFl6s57a4ghr7x28Syxnb6i3Y
CuQ0AgOq8mtDdYLBp4QjMvQsFDz1uMnucPoGI63PcHDO64vKHsKskMZkWgNedoSYhIUBCnmoWzcB
iBd7NwS6VNcsau/oyB1rUBZD7U3LZrZeeAG/hhjwzHKdYXzROp0CmNW9iRdDQi4uX4nBhU9hpc5U
IhmEOTNIqtplcP6KxDkrKet+s5fAxkb5rT2Ks1xlSCiuQDBdfuaCZqnJ6qg4TpBJOPxx9kAdpyi5
Ixb8W7mM2+YCuMWj0dZzBwpdu8tzim673+FIvSSVnF2HNMlewxak9QhfIvmfiFheOrT2yY/+9qC4
O+6FrwuPodrnlN/92HfL2wcF1buzp69Oc8snF4yNfZ3mEK8kMnt662hWO+F+YXaK5OL9ewA7whWH
jNCRSSq+YaRQS81c+tkPUujpJP1b3H81U72vU++3RohsNNq6iHFVpDQgJyr98RLIcQjg+0Px+FpI
935eHTxr5FSg47WUQ/U1BNEBhzZq5LSxoaOWbVQZ1Mh+eK8L1mcQylCS4L7N3400ay7b9oG2/loC
9DvuEyAH0yDnMZ4UGC+S4FYh08ivCRIotLJPRiFERxGjZX9WEWwK7E80FoyUqvFQJaE2gS1OvW3C
uHdyUONkXPvehqGsZyrw2uUkkmPQsHkugi4uM7AqDd9ltjPCxgIwMI4cGLrAurS6HzQ+syupvcKw
Ujgb3OZMVD/Xh4z35oOpi27np52FY0S+0p9ZrqNjWds3qgyiV8uXEEiV8vsSqZZMLXpo2JGERYzs
VwismCfdMDMbrD4JJoe88wPf044l1rYZFUlUd3LVNWRxqEw42dRVuPUe0Y9ggTC1wf6nkswX9wLp
yYM6QvTuWCD/cDZQ7rNQ/VvEuQFO+O1vO/6LcY/6xiAQTOZvM70GMai1SIph7iPQbhfivlT4zVKg
0CKgGQtpjsOhdCn5cIfACDp0hrhcgYVHxZMzzCg4N9NXZ15YijCJpo334MdtZVyOMStuqMDHkAfg
p7MuycfYEEpdUI2oyMOWziXuxWvBbjMBf+RV3SgFa3B1BdxxQuBsEO3X02dYwG0DvBeBWnfkZ+3A
oOj08sxIXHmRvHBvAzyVjI4vATPpno9Yo0YZlVMHJrTifY/8A1i3CtoiIuBeSM94nkwQ8xtx7gZC
hCsKUmVBf/O+Mua4BQkJF6Mp3BkpG3RiI1LZhuCyHc7XinaboaSHbHniPwWsbdpvr98PNaIni76/
wARcbNw5I9gI3+00Wk9RAcDp9+Jv/OPKRdaN/C10S2bD4mzJoCKOAUUtez0uvCCcy9mehnF2uCZF
X7qWJBPl22w5E9Y2YGPv69/6qX3UvgvxzlxR2ezp5tJzZxyNCE+6RN1cnuRb+8YOb8WnvncA0M5V
n+Sd80gPRcvSpWKMxZF0H6HmMByzd4uki/dZovZhBvxZKM/w9yMKjsYyPhytszDmS6LuWNAPWvu0
L4ft2vJ4Na6ckDljktcXghGgdeNkUzDejOk0W3y6mPizmENsgJFj5EBo5mIm3YDU0rRgnVxfJH2V
YRtt6iHhSQmiaOO1h+8QjpP9RMz2XfqUO2w8qoA1V/qWRn/92qnjbkljkbVlkKxW+wB1j0qQxz9t
bBGc0ewW5zoZDv/59+etQdyhBCuz1Cel7lDWYybzcmU+dQcxzitoRkBkUb3ffFj3n+8vyGUe9D5h
6HXBXK5z+i+AVoAR10JmHIjXVUZQfM2e/BLFT+jPc3Wf/Ng/r3W2W7AbditgOk89HW1hZGzSL1D6
ip5euHIzE0G6M/LSeKCAQRWnQe+S8xhbEqlqP2G5a3NrzrdgK6C4gEwDtMHC3uyqUElaJ/+FYhv4
kUOxcxnKHktyvChIgI/nYhvz72x0ayuTRUODo8QkznzVsdxcboMhMCgb1SVB0Pb7vA6I/lInxxxt
D9A16koobfejEi9RJcEdkmNqkXQMx0ShDkj3OrDYGKRvm0YEOQeVr/By+QCGTRUoB5t/+WHEa3i/
zz80AFQdzVWxnBlK0AIWulG6LRHcQC83h28ehXlxmeHmOkyAybZYnsrH8N9QWsDXXN9hJVqRu9oN
bL3UdWSDZnd8fB3Xg9eIf69qpU8vResRQwqa2KE8P03c7gL/7xGHdu7UE+viQ5Ki6ddBB/K7mkYs
705XYQuC3JkVa2emyJIFH8dmV1xoCBa54O9OK7X2AIqs42HCFDDEJ6RwTyFvHkHVPtQFq4NaEtGu
EzNyNToALTbJwMeOIu0X0u60S/LTq2IZYo4A/hYlveOzq91NFoGLGjs+5hgAbWfka+RLt9bPrAf7
A+njvFthMdgUCz5CCQCvnGB+dHhqk5B+hi5S1Q21Cus1dZzPrBvpIhY8ONi/BH3j3LRqYnxdgNEC
XSZv2uwGAVPLsbUN6DwxQEISZ9p8QBefamqaKPDJT5pTuDg2HANQirM22dqigmxq7PipKa4CDyrW
5/vA52f33ui0uTCmyck4EFdJ4gp5V/N1yIVIYEZJr2suBhDzWd5zoO3gJqlmq/ifUaT8QsID4H9p
/omBMPChUq9L42C6pvI7DpkEd+4RmZHH8wFhbmXkjjFOTxxOl5rB0wdBtz4WK7Ro8eSuBmLdlFvP
tUQBqBxSPsfvSd8AB7BTF9T6AT5zfbOz7Xp+I2v9erWFrIrjDqjTTIUUvuii9vLKnG3C367hAhyS
zJlq+jgqnSAwAPjfWQ+5No6QNE4W4TAUAlUAVeU2nC2xSOy99EJpM6YbdW3TzW/6DNn6YrBlPP6p
x84xgL+nZsInvESrreC/yCwlsAE62Zd3Vah2Z9gXlwbtk9PhEX4gBej5wsLX3nIDgeY3ZlRi+ATi
94T2vuq+oOvsosGL0H+cY7RyhCkwQk4SI9EO44dHjIBtHINB+uX0U/BwJyyiRLVORxECveAuEXhN
9mBCqaE27GzMV9/CPalqyZGchVjAif1+xEw+ZeqyfjEVc7tDIxAB/bo5DsVSmDqVs4Axw3YD7E5U
qYf9wYhixECl0QGfhb9vdBJzjPG2NUid9G71a28prY2esiX/LMQb1ww8HZp38Y2qGexoIQl2m4v7
UoZ+ZYXXrtn/6CXg1fKmYy25S8qwU4XoTOv6bmCEWyhDisI6qJTpI4NBnLR2Q2lgGl+SOX0RgamR
D1KAH010z4POhuUNfnvMTijkY8hGMR3+E+oLEweeZQYQjKi0eFlNqoJJ3kgQXPyQ2JpThjYHBcyE
bYo7V+PwRDh8JzPYNGNTPZ6K2Z9n/ZppperL8sMVL6VzkSPaNmsTGdotS1r/cHnYGundc2eaVYvp
EFULS8Pcs3gQrCouX9kd7L5aY8g9pS/rdaHzSvOMzWj+474jFJQnMjnUsuW5lbz6P1IOkdi+SEZS
hcZgyT4cWuOmTD0TK65IGfcie/hmiDpQDGsPyN3iQN9FQVoEK8MEPC7UmIdk4Pj/7Q10/TPss2wK
w/9yOX7Oc/QbmOWDTLNzSYNMvQYv5t8Ia9LJm+YmSz9+tlsqZnEr0fPUIyV92yQK0kiot5Ne6tlJ
di0kKRQVSTm5OH/5RiMd1pf1EpXHy7chn9o/PfrQxSvTw+ODWEN2BvFrCCe/V4OOVbLVeLbm/jOK
cMH3gPDfwU/ZgtpGpim9jXcgERhAlluDwQouo1PvBfWeUuMoQIXpC1o33x6FpfAmdZ9nGjB6Z/3g
OOD2EjeubJpJA/hfMRe8GmncqzlN83jWzT6DV4PtDmoARHA8CZ8LT+siJC/yWQk70uN6oBjWLfaJ
OfQIxhp+dsSrx16CJd7MBoOG9RJngaFeVreKfrtJOC/I1Wd1x7+AOjScUFA5g2DFMeX2POvxkRr2
t9/t3De57LHNNVGvPS62t/wD78a1aSC1ZZraw7G6cfs/BgHWraWUvhY+o27WvpT8h4A8GgPCF8is
kaiERsdZPNvn5xu3F5/BXRQaKW4xj/TXT6L6EfeOwNSDA8x4Bw/+tslcn3FyugiPSD6X4j8aEZqR
2snfxMoyP5ydZ4Ab4L3EFJzRFG8tM4oAvq9l+buhB6IbLV/9lHevENBH6BGOq6zeIi0PkPoh3wnS
G8IVwE8j8eFwZBDnPozNQoEzlhOuZic8eN0BF7umkCP5A2Vqm6bdF5UCWUnhsdkRT5ANnhDJGOCR
HWUohT4pTcqE1S6PgtFqk9m4u7fo+ekIMBJvhi7rrPfAiHaGNirmwsgdLS3p5FnZfEoCLY/tj4+f
uLiH+3E5ddWGX5qKS9xkeo/HT35Cl2PwpCq9J3wl0/b+IZDc6tbSuLWX7pG76rzscipCHVXBzYP7
AgjX6lqCiB3l/QF3UBNEPKsKUJaiG0R99ax9bEiKrf2zlQfgXi/tC3zspaYkKY4U8Cw3qxHiLmg/
1JnWuXA5h4JpbKWCl5KoFBzAetN9XmFk2vrM7xdAs66wUmB4jOR/cUt9GEBvktIc8f1zB9AC+c2S
52DbvszSmD41FEgmwn5XmTuboeqqM6EUibXM+sP6MQ2TQkCq94iONS/w7n9nYuqRovr8HOkIYZDQ
QU47PZp4hYQ4Qo8ACtZHcjpYoDNHKNGAGCDpeXIcVB0MBua8qYUUVhxVzPLb5kb1wbtBLvc3Iyfi
2fnYY23HWjBRwwc3gklKHlzjUODJiizEVhOKV3Jx1sEUhpoeALvis/RuGYNdukkJD/D57LBL/67f
q/WPqbGu5VXiMe4ATNi9J+uQ1xYUdIMFYJctaG68kOAuPaFOXAAF70tqRp62kylo0Gv456T9r99o
Hy7kE3+zAxIBJ/jnxYCN+nSJVJlm1U31Zc6389YpHOI713jzLD/cVQ68R8ST7aT2oiVlApNKlwaz
X1aJN40ub/PtyI++90PiP/Gl+MIUvaDPXq4G8tVPoDywzb3BX+FUm37ZRlDWCytjFyVOK09+Cf9p
O/EMIUKKxOTYcx5qEQZc9JDGHU1VKUDXVuh/vcUSIuR2mGDbO3PDNB8+vs4Z3rqIJ/k96ZZlmPx0
srz8/un2l/N3E1McQuuVP6nVct4hvf8X+Ts1dJMxRD9MVGEq7IxHGaNt5UQssFtce574p6RyMIdU
AMbHKNnt8/ojghwZ+JuimTAgSzsUzTFGDLiYcegaJuDcYmWoqg+bGFt3ODyd8RgqQnpoT8rlHs0E
LtIFiXn+zkddKvCJXSnb3lEbVN5xPAXu7elalFofhv01s/mHKzQEUAjy5oQlLQruElQSN1pa1d60
ZwuqMR8l9bo5LnPFkAPab8Ft8Cqlkw1e8j8a0bdiy7JjnmFeIKJRgBKxBzwsG/AZMtYYlzwmg3jj
Co+BJWFa4beeimfSPOCfLEBc4H44X2mCEW0B/chiPEcQENHxJ9ppODIRn4GqFdBW9YpSpkTtEIrP
WoY5W9xVsQ0RQc+ErOBzSKlRQP/j6aXzND69PBjEZgIaMD2OXlTiQ2tpleYRwzZ/GahVy3c0enLY
szo3wqkvLNqLt+O6KU3QXfvE4FWqlZjdi4t+2AAwIZdbUtsz8vqL2Llilmpavo3rrGAdY74+y+av
gLU+66CZTwMUPNfsSW8n9WN6+wDjUsqxyf1yWG0Y9N28HVjFPrMZ7O0MfGzAILoxYH9a7x9BRAdF
keK87k0Ubg+Y/tKwPKapieADukvc8C6sfMKqOfRMPhUwOfeyLW0k191NOMBZeeywIHytEa8wVa56
H34JX6alY6fGECTypnhpPHQ/HncY+WQGkrqu4EmPa+HZOamRJJzSg3M5/9RxPCyvVUPb46tmmjmG
9KD777n4RbXD4GhUlr1PqzEuvv66BbdX5uIvp2THBe+vV1PKNwUl1CGVJQIj06q9oG0KtOIrrCxC
A2KUMwygmwxW4eMAb0MIfLwOaI0qTnGeFErsLghc4XUohVzjdItMMrsITv00iX7y2afZxBFii+cB
HICSpQWXi2VWNcLQUyYQkiCc6d/WdgsFUbFiO0qOQ2N4FMyQ2GdodfGHmHdSM8ZLugG390MkOiyP
UEnmxUGXAUcyYQq3OYjrMy/ED8ratc0dgXkOQzO+S3XfLlm7lHRFw6YgWz3/N6fVTKdrRpI3R/tx
gakqB1YPaRzKLz3IOzehPglXI2M3r2wn9CyylLcDD0wyk3TpIiCjuzkdc04FpAHXsz/D7995Yrij
JXpIZtk5zzmPQswYxvRszK9RMuY2Ajl63Kq5/vTdsLXd+War3lJUr02E/Gv044JpYg6YPAiT8JXu
bP0UmFOq6lrofDunhd30RZAGjNEz+U175yfq7srU6TzE8PWWQu+MPcOtosrmmdBZh5ALgcJNmsbC
qcVzikngsUWZUeNn2IKf72Gl6+ndFnfHCNZxdJrO1XiKJmFBSZBPJbm5S2XmR6/6zv6q8qMiDs05
mLJE+HqJtU/V2nhWSW+VNMc6O4+vRkH7R9P4IMhWR33DfaRoCTw/Vn83n0hScMb5R0BaY6vq5658
G4x8nYLdkk2qKcz55XqE0VB8LTsG8ptAmIx0LE2VzWAcxd8tZzoRebo2kuqWrhr0smJUWPnF5qvd
D2w/LdqBqxp1oKa9MgfmvYmvwEF8SfG0Nt7lyJLCGPyJZ+8mMWqB2s5DgAXfghmGKHLzeFVbsi9D
9Caa0Kgrp7eSKIoxNWRQRpXD99OKArXXq4/H1T0wxdEir+CkWBik8EFG9sUhhJshhfbUxxQjBoNQ
FGX//J/uJYTobaCS2FZoz16CAYr9m1MDOfvVJIvs4zU9HyPa1MLDIonwD/zeC6mIllxtAc5ZZbF1
QXei6af2LhE7VcP4AvMRnddkkAtegckqXUzjkFWKd2zWkGiS+hsbZeooTie07g0DIkmv5L04Kye+
UW32YFIruy5IEolahoWUv6g+91+Pz8eZcuhYYynhHutCYIkPF0y2MLtnpToennvveiPO86Y0vPYf
wJwsr+BLD2Z84cOdWgyz8WTC/TMGxNcbcpWvtFEmXhscf91ACBdQSFBUclHLUGtnUKZfDGpDqfqL
VAZgs3ajRrkdLrsWwMlMn3K2XeqCucKwFfOoM5IzVksWzXjxb9onh2MYZGyLE5wESHk2DlzlI+mQ
IttzCmeZ9K+hQVguFAU+qxI42lcJM0qE6uqBcZElwexq70fkcAJL/dkxZoLpQ5WP/9zIUq/MeIiS
iqHWewHp1uQbJCoeEkFl0kRxK9eWF3z8T85WSfIgdo+5pQIw6+HzBBf5wbm96mrG+yTdoSBgsZr4
9ILLCfvLp5tZtOtivOatrtIQ3bPGzczLcWtAeHRuEdAxaqy4EeS9z528Zi2qhkz625UufQFvoK1X
/j7JDat4J1o0oToXHhz2fHEJoE/CtwgH1dyEKayoqcCPya/nh8vtrkUhPTkOg0z+YBomu0o2zZoV
1sOQnv3cpQsyu2LIR4KgQvsW0NbxyyxCpF65Eu5ifdSdo4uk+nwqB9oTq+rdgG/HhEUvlk/4YrUd
e6ohVBLlrR+XOL1eXTGEwLFnVdRu0/hg5PkS8CT2D7O/HGD6HBxbFZSqR41yOMgJxiAlTagzZ2cE
87IHu+e14E6E1Mz8Ux+t9VavZx3eG+rBunncaypV4JrXFw1gwR27vhfJxinZgZYRGOmuMOR1AjNd
wQvyHunXtDsNcT8A5ZTolRMHGBXp/gUcVt+sxVktPTn5kGOa5uhBcHHi1Y8eoHhlvP3gvM70Ql5n
7ebLkFmEj8+46Qn9NRiQlAyiWmwTGlZNUiepppehRdMue2FNHnzzxnCFH2BHZYO+J+PYlaTyQwqP
5enlPdGE/VcJgnygbB9PiZRtq2ceYdM/ADezR3U4yR3Y4AqOuvI7GdKywlwA/qmzY23SEZhAI1fu
/zF1Zkz+Yi+KQ7nGUhhrqzSH8x565RuE8mS16uKU++qyOpaHfxWnbLKARcI2G+QlS0MHqzBtAPXP
6EmTXE+EmqYMwsFnFLqz9q9dodfkyzxlzvATi6uNe3bkQ/ZVkzmoe5gR90kRsTurk6O/W4hdoa/o
t0xmJEAQcgjXnG9Ux4m3VUzVPDT0k77mxnpO9hj7lZIyCqWOyG7sF2GqAZ9E+5ucx31JN0pWvrZQ
tGhyx0EsKHZB0NHWMLCalxunSQVT8GPKGTmb82/cWgZEJq3TB0C27GzvwSyQGPpx1LgAYxTmO4u1
XVS2Vr4DVCABcyE5Z5zoIVfDPFkNlpD8q7z38GLFK/LWbHt6MYXLfycwKEOHCvFWL4hTsODZDrjn
KA7S0TrQF2cSxVMVmamIBh6tTqedMgrFPQzryL1bJsO7xlsnUXqsKHWMTt7Yfy8u05KavWGZq1Db
xPcP6c5jamSSb1zeRO8duFzE7QyHHq+EMJ76tLkFSmpT6Ir1SsYhpMbqCwWHO1s5F6Fy28BNU+4m
oV74/2oyfUgJH2gajPjWAtsrUYj4NuIFJ6WUQanWSqfmsaHJ9B2LPo7kXFQkDy9HHUkmSzjw64dV
aaOOSFFThWpfXm+TP20Q1QbBefzkP+YiqbpHXjUjlYmfuzWrGAAUbs5jl5JT1uh9/m5yO7f1zixp
QYb8zgQiuOPxVk0F206MNdjnCPCWzypfF/gZwPweaqeZ/YcOO3Ue1xsclrKEOhpabS0dPxeexvUD
NK53ad8VowoMfJYqo144BZizXztzQWsvyvG7Y068s1TmipkMT1bS8oiB4+idql5nDmv1devgv+XL
Tlb7l730cMKsjazD5UlY9+6GlWqKhl5U3xPsljq3yHuN23aV4dc2J0p2vdi3iMAVC9TeQ/2CBISx
ouhLo1O4StdJz6uMav3Ut7Q2pstGHMfNynum23RIboSrj927pFPQ2GQXP0xjSjcybajspOwwwsJ4
zNhtGS6Hd+V4IwaTuXCHZnRV/BL5GY6BH+E/6cYOk72Ohpcst3wwiSfnm/I3+ndCkQbM9+GJO3w1
xh1jNFkZ8aoBs48fDPnyTxF+sXlxcvXbV3bkHz7rkGvADQSYaXkKVik/KxtMZ+WDmXiK/ZP/1SVl
Xv1+qEH7R8EfPhUaDYRoUsznLJmWGX+bwyg6Wo6CqW4W8lNTm3Ycvq1n3WoaLlUIfs6cv4V/RE4X
L9CgT6SKfNC3ez/+VJCfEF6EM5NmiFi30ERziPnr6q1KSysZBH9qrPp26Noc9Pj9L/FIgxvT/Xdx
lt1k7bfDhTyWDX3oKMIXl+LGU8AnJ16UsPKP2J3H4rkGOrfXCC1idtMuFsZyrQCJrWARG7ZE9qUX
L7+kFmiwGvioywtvnanTQ8vXepYlcHuzeGqYgWMDMhSlwyIJpoMr5gUv3utpqqoGafFIbFjLgAVy
Re/MXvVfuQd+Omi0zPsStS+wjSYhkLlPwyVYxnXVkgGu8eYFrFK6NAMC3q1BVnQ7tA5A1Srn8L6n
TbxNJ4efG5dgghE0QDW6w8K8/bZ50bW65A73bk2q49aYPkZZ18Z4x8QzgCXffr9eVI3O55Tglg1x
iIfw2KjRUO0yq94vm/s+4Z3q7JKglgWopwSpV9aiVepsxh3VrlWus9/DpKa4B3hOtPr7g0gn7ewP
tjY8KaUUc03LAgGXKCOkep2BIMWIe39/+UtB1M3qNEiQNv92wvQt78tCOS14w6k3lmpR0Sx1mjgD
efF8VFDmfnNcWPgHD+++aIgBnN3jcGBey57IFgiuMO5qigQwbJUMsmTkpEXjNr1jT9+X07bqzgNW
SzPXDIPckKTYHmtVE4DACFVNgjDP+Em8ScWKrgPw9ptrlDyOdgSJYxZ9e4Dkadz5cpBWfkBuvhzB
P62U65tyG5BmiJ4hredpPA4f+Qs8A8qmqxYwH//Wju94ZW6xIeA+H1u8RkzmihzwOpXsnfVrIcEm
/TaMRi9buxfyZEQK1/t/kXzfzvQxsyhN2pbOB9HxA03gQ1MJfAAXhatxotjb7d0rs5UBzj33kTps
2qmWh3Bh39BgBxHZcNJyNSb0cV8GG3oT21sgvlghsneGjMd5LjkzhxDJLWGJQCOcJFytN8nttxkr
tZ+m1mAb0/Kb+rrDLfSXl68fBiGPNTYdK3McYptI+NfbaiKvKzZ8wsS/LPC0yzYELtry2RlwEhzF
62PLBmr7vLPzSJcQPhJf6UnBtLm6+XJFdtXjWzLVFYyaKv76t7GpdnJEODGewbSGEUArNUJ36ZAn
uv23aFrY2PvFW6toCStoOdLSI/AsXl7Mt8JI5nPuEbThvgtAhGsPcnOS1Zjch+3sCTmTERQvbvZR
zyFBNjTJw2fQuiSGwIwwIy7obaL2H9O5zCmo35iU66QQAwihzcSgz8+r9IU0ezwhD1SgjDRRxDfc
IEOtqAeGlXQrT+c+7zUGfYu6uAXrymhXygprAVAfGrBWwmu5Z6oUL9WOAxuni6FDiesG9jVvjocd
pbBCwKhRVXZ5ohmoZoH+QBfiJxf/mf0ifRhhLrzYEKpwwTjM0HO2u7kVbhsNQJzTWZPpqnsHsuZo
G1dJ6ufvNgBa3hXTYv35nnOTbJcQ3scJpHZksL1LtlfC+61VG5urJ+Bp8Rc7HScR9IE/BY4xVzXw
rVTMquiuVNWcDNQAHYpZ7j+vNiAEomGUvXamB3sKdhis3FRHTiPddIjXRO7RCttmi+AVrCVIEHXG
T6lv6JPU2Esk7zzkHJr94pm/ff0KgzwWmHVv+57cgOdu3XeGgVOxOl2Ej3vwDcSGQzZC4wMrubNk
B2y2H1frytJu7evXP3iBhxRRPsZY6gAuzg7SvhDRFCxM1Sg9emONac90Ds+LnbOMT1SHNEaFiqH0
nPDWqP+BoMpxRr+7eW3os/UclTCxCFw8z0oPT/eqTz9s9915qV/+4OW5jVA5RWL1grWtovEAzXCj
f8m1L7kx4VaXrpzdwMUIAvRbbH2i5BLxrcv4o3B0lmZdkgd+Znqm8ThbKonx4oDhKjTKmAS6vKVJ
+yVz14n1NjrdHyLFQEz3AlaP4rOZhAKvNEBGyWtosw1E5zb9a9jaIhDQnLyyOVnC+RNtDK4SODJI
nqW3HSr91be/qAnCEzd2hbOLvMvIYyyR62wSyJrkO0LIxR5hMa7FCKrc8xkPUkP5MXmKGN1u2usA
0Hi9is6XiOyix2fwY2URDy0xxi43ld9wgd49ytqAupRTi8kjI53X4RyXUPNUw1KCXY8I3a31yQ8Y
l6qD4cIEMhLB+PrRAlHyoA4l2Uy/CABH7GwCafYXei+3fZ6hABGFLA51gVMl9t+zzHiwsgKOsVMG
tVjkg6BxXToRxa/7+fwutg90hXJSrT0HnUJbIx+EUXAwkD0TfmhBothlQ+OL48lK++QWRU+++BSd
0cLlYz7XyI4QguLPAMTo2n88sdrArBONzizz9talmrr3jukRg6mvc98iQ30OtrhmCPCqiQTLbcYI
qip6MOtb2VWP/GRkeBJUqoSZZ9LJCUzAnnHGKV8nT6VnnZX6VO+bcTsPq2HJk+vTKNv+rBWDHIv8
JN7LtS1CEMnjs3Cp4EZka/Yi5g59NQvFzSn8UX8MUHaold2bmwDtn/Ll5X0OPNkcKxCEA2IVf5bc
hQ4CqHIT2LaLrtgEoMdpTENMSC3K7nB9f65YmmdxHIRcz/fM4elp/WneZFtGepjts2WDN2ZNwawx
TBB2cn4X5ckFEryaBFViRUwrFYtAxVtpaE0rz96bkfT0QoSPPLelVpFIPioSGfaVmsGLbvAa6SJV
NMddO5G9GjEUoPsBbP38/NdM0OAkmDWIqZK3tiQP6Q3PZ2i8ABgZcLIA7LTokMnS5zMYQDNYD2dn
0EDAgyU0bPZcqZ6pbhIY2t1ERxlT5etQUkN+cfdVQo0hSY2lXBb/GO6/zhj6vAGFJgZVIL5wUhdb
vnMJs/LgxUKKNQfyOiVvc5etadbrL5yJnPnT0NTKpVNbO67uhJ7F87rSz789kB2Et6vuNnwqMAek
43lnQYZdPisVCZbu1UImfhDRCMIlaq6klpbBotjrctc9mnZut7HSpc8qYDVuqM2mVYlcrP0rNt5s
0vDKWAC1XmKyvX/rBJJZZ+/nBZrl++xkqMPknGnD60SzmEtz1rfhZOuSGlVtmI4s+GfRATyvRqgs
Yzo+9iGNr+CyWwtQlqTuFxnrSuVlups4WpXFk0X2lmGJjTuO7guPvJFMIoncBkU4VqLv98D8mAiR
t3/quDr21E+WTiYgxuygRjKcItZ6vTgF7GMaS5tO/O9qSdyIDeqQmz1N+PTYCzbiBopn/1IkejBV
jeVLYkpRhweeLvP1/jA3IW0BD8vJPS4uhLa5a1A1BWqBn0z0xk6XBSms8UgmkZTGGEQKaT1SGkxr
mSRIr6nB8ugX5lrpvUWLT2pjcRYVeTV3r2BW+TJpLLHbAtD7JukYUFzny+sZEWVLvWPAFZxcpL4S
v9NvnZHggONKaV2TUiW3s++OU5KIwtyq8XKaIxVLjcxtnvtlS51gEb5y8RQuDaW1EnhiVx71tXx+
GqVpms/wNHGfhHhn+qlM2YGI3al52TujN4egWd+gWJrYuuB4bu1+zKQe0B+LwMCU4Mgn41CXmCGI
0c/T84Gas12dT87TvycaiYUn7wWGy7FnDiBN+RfPt88fXhD1RFK77Br21iRugBFkxWxb7mvLe0g9
apefVjephxte4+bPFc33f6P+4x9g58teAFOw405SJwm8NHxc83CFJkIu6OVzAEL8mRo4JbNwQfBe
TLCUGtW5UvGkXNDsspEy+x20e6dQh2H2VZeAj3FRdofKjIqm731dUxBXXlGRGbGLE1G70zH+c5QW
CxogvB2V8o3YZ8Vq4gmLLnRsFEnKJt+FyVqVDSds5zoHIcaYFrDf1aL4iY3S1FtjTa0JvWZ2UWgV
+9xajk6GT2O4Ox+uhS4/zyzjuE/IC2R7HbjnTWa8AR8NoCOhcMhl5Gcg/NJ3adl3m/vyV8M28l0Y
OWK4uC3tRdDAn3DQIeg1/dtF5swDticRmSww7N1ifn78vP8YyfSSGqEpq77dcQTxkxOqd7FxYMUR
vfwKHhMAZSvCYxSoFBo+ls3CyS/0ox6X/tb4Wq82t3TIfUnh1CaqJKZcj2LMQVabV4ldkr5XiOK/
gl971PzrZj5SBEaMlstS7HPKB682MwXU762cCuQiZJ7K7Y0ng6xOasOAHcAsKZO6GLAAUwZS7zSZ
sWIieTaUCGBuASBWbdHimQPx9CjqlnE8Lf+s/jETK7xYP8+O2D6p8cvHx7OZM4Rcn/CXXWWKTAkr
0/iUShpaY7oQyQrdSCiO6tzYgJ8wW+jxXBzMjMcshk02krZglk1m3GSvlxERnuft6RfYTVncPSxB
TgXOcCXrlKsmy2vnb0Ei3rF+0kBXKrZ27JO4deLLn8QBKm3O+pV1IabXOR6Ksh/MnSakFCOAnr2o
MnCkojRyF1W/RI/gtKnJG+Twjt8CmCLZYsWE6nQCTREqa4LKyVffTCGPETqf+mxJSaFR8Lpt7SFZ
Ew4JrW0iussEI3GGsQsp2ccTM9ASgf68svHcUpb081Zz59/yKSEyNnOPHApHb8BZmiYHJa4v/mwy
EHPK4y8w6y+o7QP93O01T/zbcUcVItg9+VmzrbzOJNtrQNg1Da/iWbH9rGwnzxykzr7nWPivzEsL
rd/ReTmMOg7rGiWNKggOsCCYb1LCtQCn2aFwKd2v14IxAQpXw6akwGqstEh5NpwAk3VOg+vsbbCr
3fW7sh7LGMo8q9Oo6U1DiWCem7OOYdSltG6kkThwKMvHHemQuhRadGr/9yHLOnb4BcMtUTc7Rv1+
mCXx+75LpxMpH6qOTwPchqdJljQXTheCRcID2NlfAQLLA00ro65TidbWJAx8TKSUwl+BXCXHBQMT
Uya5SFrvyrgj1kEn2b+Zhi/8KWeEodAtJwrv4AStiLWxTqjBX+eS14O/tQoBqkkXU0vKkaxVVleI
UPMiHVnjUMSWh4pQhOO0jf41hmDLUAIn0uhQi7Hdm+xUwIAJKM/39bx/wOFYxjjEMcpXwDdbk7G1
yi/YLOmnuUuodBkq0R5diDw/K45P/kg6NmE2D0KyVvvlWznpbYY/tWWeCIT83YElvOnJg9GbKnb6
ZLF42+Hub5CjSakdfPjT+2Edso03va4Ub+HYb7NsS9qMnDZ9bGwKUgX4mayaTEBqvpkP6jtUo16M
/wJ4QeyrplEoMHUdoiyjiuf71yHdgFV8pFRUCcYQUPdrDr/Ec2SSMsT0jz2hVh7EQB9U2aatu4me
+YLjUQLEryCWnYl+tZnPmgGcNtQA9yh0tjxoGU0P6+V0fMk3e1wcnMwHsl5JdUlVWGwzGKOFkk/W
xfODvrN9MK3FrjsNAeeNbz+nI0uB96iy8kjtBJMOCybjLi7jLDBNrYsk7cmKhqhUvs6K4tECUPD3
5BdXWjilZAgNPMibmcyNK6kx5w8uC2k0CkBewANHX+iAvVQK3nnRYpV2xKBiSjrN3TfVXY1DISYI
2BqV7sSvVVxMJSaSAZM+6O9O/Uoq6Y6s0K3p8FGUYkOW1kw3Rx44aAwvKWMcUDM3ISVrCrnglVRV
Pneum4hP4VODaztlacLw0Qpfz3kObRdktguZN5bD9wXoZvr7EFNXYkaK2PbCSpPEr8hEmJCj3PAZ
Xh/vcKLIg5rnQ35HadZzIpuero8rfXpVkoSwD8ZnbNsGjjmXGMiwoyVuGVhUl68zOkjP77MQRKB7
USmBvDU9W7f0wxjWIfjoyoOm2BgQyowkcUwtA6SjFkrUl7G5+dOnbTXcCPnwc1vDPWBE8effDoVc
8O3gCdvURtffOO76j/IY7suj+fyFGL7rnb3/p5gPfS4ZiKiELQw+lA6mvX50Qgk4D7i1fmBwa3u5
ELAFFVTppNNQY7F1UJkIxeyMCypipBR5TEtxdvg9Qxg+770mwk9ZdyQzpezFfkT6fMpAIM2T0dZX
6aEycthr3zmVJNBWA+Xp8OxfSo7SPyY6SfSG2Efotw5o2Uvww9o56ZIHyUbWsDuV+Vgil53fKvWn
HNwIUm6Job2bx/3Fm9FEQ8s6ce4W2vDL3TtsVD0DsPCV/tm7X/dNpABmXiuE0mM5R/6+JbHOjP1y
eOOJP1fb1NAJggitA24nkSZ55ek9e7zCkI/uQHJObn7MLSkQBAmepbVgODT0jpV/ShsVTi1JBGE/
eLT/Nj5xzODAECjwy+z7wYkytnBPm3QLclw4UMGWXnAmHBbwOcaLV+jLroYwvGBsKx0MZprx5uQj
SCKtet+xSQcZB0ccOohdapblxtrSb9z13dO6J55TCaHLcC0g3bIprOIe7TsrAW5Ad5M+qVhoGPmF
sjK3CWEaGuODpBo8r7bxeG81vIxg+nxSmFTmtWW0VgTWVn0U85VXRCoblLDxvSGnP5/mcOqh0aq9
GBFeU+CYA7KjQuiZuN49a2Yhmcya/vLYdy5BmIg2EfuxWzp81KmdeMf6JZbXJFcsXoedSoGikB5h
BzLzZBIvW/F6tTqPMURXO2Oy0SeJBm5+JXJiAFKkf1PYMRqxteaL06yPv7d72XKoo5LmtYJMzCvF
JitNQKazNZwcAo5kVnZqRViQlGwwl0Fp4QQHdLQXqazWS5f94kU5G2VjiV/2wGiBQ6COSjT357gC
UkMx0RuTvzNMGS6+uNSTECOLkxAUILSC89X7in8/IJ1GIcIWa6nQZCoXUPCTKzOt69dUQ6nFDVVM
HUPI9hfUtM5hFwK47/OiPl4ypNtZUWyESt55RJJJfuLArKSjVIPxOT1pWWYhUtEVgCyuLoGrnu7e
Krq2XakAgwTjHnM/TPH2bzygVfBTPpOmbS4bbyb0zBD8RdtysjOnWayfdSwVI28vb5CxOcxaYjS+
we06s48WfpTTfmhqSYJ6qY2Nc4OXG5mSzkjCVscB5AvqCUBs0KY/V4yOEmBzIDhr6br2fEBytLxu
SzwWev3qwzOG3iwOORkZTh9DO7TMI8S/EwcfXzQzPTJHLut6thOGukjet+cdRaoqfJELfEEHEsml
zjHmONQHC+lMPsmkF3/Bf9vtNCh/MJMw2p92zy7oQkV7VXpOK43vwxjYOPrn+G7vTrXUt3fFxVVe
uu42ZTnH4u+GD7s2JHp6/g3nO+ep0FDZRbF9v9F6aZ9EdnZQqTOkpa3h82c4UIet1wS4TSH78N9+
fH/zo8X8K+vPNsmXIEXetswWAFcPgDEwPM1IhQWCkWSyVPNmi8X2D1MQOWq3TEMWsLm0BAU3l7Qd
Qhw3zHSoofRSmY+PcFE4f20u6dmdUUnVYpp82dMwtUBArLmBySOTV/cytDyBQgIGk78c/779zRVg
Jzli/UVxls/bqJOR+b26mjT0sWeWBiOph/MlA7Ikgw7tZHABxbz+fGQDhIzV+HxQiCAUZHEXQLXq
3KnBKmi9DZf71+tw7Oe+IS2OT0tk4/au2t+S/QUWpbJnLZG+peZDpdYaQclmUvK8RcXzdvGh39jj
5FcjtaKJv9DHRnYtT1dBSdInG+cRKEmhKN3UujvGj5+x+7ocDgaW33mubRYH2Kpplc18GYGL07bh
lVhl6bbEZalXYuWAkAxlbXKIS1j/zWGobhEspfKprXnEBSkr5uJP1tVH6x7k4N77fC3bv1tiSqBG
sHlGi2hyQXiRTYwBdQY312H53CMb/WU23hBYVz+1BMXQzlaPp4LkHg6y2EgAXAPw1Xzj3ynu0xJo
f4lk4NfAgM1n7C7b2SmEGvK4o5p74gVg9HeQQGIYGL/tSb4SIPFzIhdx8C0B8/sdbivrq3j0SEJm
uCv8lTRJO0stAgMMz27glTVhxwBlfZNwi6cxCivGL6JKJzYE3kyyHhFms12zLZj/r8bzvnihlgVo
hoJuqX7EZHWdzQzXWEDRY7tWXBfefXGul61PjgHw6hgAkgHDE5ICgGsxLGmLufiYXAEQtczm5vOd
f9hGL5AmhEwJE2FCD/MT+NYzU53JZ4rOATIUg7VvrmB7TvLUQzndTCmMf+eLVYcRVq+eoVwGxrkO
L9iozQHMegozNZa7e2I4/bL4Re4UbLxFlrEE6k5iJQMT1afbXRs5IWEHcv968Jy2584Mc7ji8tiB
rPx0c/c4YxLrJiLM4ImSNKIVnOhSNn3+dMu1aUj8/hhLhLEy27ozycHwAfHQdHp+XMEdgSrDlEKU
gkTbBmAdlVNgeKfvWc6vC9XRM1iWp5XTcQMrV3MgB00sTNwubDhyuVPNgDNiBjbR+bDIKIVaFe4j
64+lMVOpXFo8nSSUhitbxB3aER/710ClnFNvdba8jN19MlQoc/PuPQfCYQOy0jmWNpqvFmr55dkg
iTmNJwvH/rtkQkPZYKYtFo6S3mSzYYV6z2tRsUpwWUqcuZYRKi2iKQZzkW6nAjO9VRNg6MJui83S
xOwrVzodrXG5csp5yH+LP6zQCkLBvrXSOUEzfn1G36gPuwrRXLGWCgP6lnNOq0j7PjVHUP3dUmla
XF1CS5+zX2iCaoMLEIHw1MY9CAPeU8d7I9VGm/VODm6yuyuTfIkN8p7q8U3PkRs4SC5B4kbGjR7b
Vg4VyFD8kkekc41fhYPvLM8a53cHmi+LERZj2Eotyi2p5nVs9plUIXmPuRIl+MzE0XjO0JoXqZmU
NXnWEhyKOsGmwjL5Gd8WeKOZn/2qplKKcJl2iveDVQsxeLAP/UtT3GrHds/ecTnVX0zpZHCiCCcG
m8MhNofpIpL6ONOWVc41a+6pAjh0bKWhpCx10lHvrvpoXF1nAHH9X8A/ql/a0RWCKFTcphJKhWj7
ns3OYA8FluHsEtLEL2DvLKVyZ+Ys07ZrFOWLt7CFAcSFs8EaXTvtpV38g9GgcbLgXsUDzlK7sTKg
zcnQZc7UPC0diuiPQQ1AWqL5Te3gjPV5SLA25zX9T5tOEln4FGJVoth5iXJNvG4sM4vDsz75XaeE
bvJlC+i5r7gh6xhe91I9LJ6eI3dUNI9Vrcfqz+cmLTGgXPUy6F8mA8bUh63tfjXj6apHU/LA+djJ
azbk7MrFNle2pXiiQcv+SaR/WBxn8TJNmBOU36R4/b+iLZBfSxb8es3ofuGyxVlhiE5mqmLqtBV8
usmEHgw+4+/cuRWcX+yRHb28Gh5vqmGFjOcmaJmy+Ltla+9l+C03Asv6TyemycvCXmQ8v9ZiyYa9
wRo8p3lzdu7A98c+l1Ovg+HZ844Elu9oxBSiYi05AN1EFD66wI7arCI7Er+aJAxn6kO1tZYA/E6o
k1YkOygsh7MV4mHUF0c7XfW5uTaB7ckyhEzLTbp3EUnvqGgZYt59EUWRQlYrrG+Cn51K09VitiCB
iVm/7RUFrll/3uNVkMKdSB5VJ8DbwcHcRgLonfIgDN+ofce9U+jsUCQaGTOA85POh25dB5nD1Bul
flXyjgoa4pI2kwkznNyF30Ks8uy8udotQz3M4sgYX8/FomgL7boKEBbiyDaxOhPJnsyZV1kp0/S2
bwSMQVkDhByi3pGa9+N9/6XhjBNsRpxjLREklGJh6VEWpeQ9a8/IsU5LhmWwvsyRsKo6FzyDbBxj
CFnVqrh7zvGO/f7bv1zjucE2EzhnY+VKmA5HcgyTarWUZd0f3tDECAe7xO2v7MV8JBK3ZE9RzLQA
H8yW/9kq4VwdLvPDCCc0Ego8pRpJu1hsFHo7MDBP8rxN7Na08gGhngjXPyJPlxcRqq5Kr5HIfjTu
pmwtgeY6nNYGZ056jB5apdCfhqhp+k791oNJH+NuGrEsNnw/vIeWpgTN5sTmHhqPH45azPlHd8Br
uR086B6Li1VbMApxeUjrPkSZUPAk6crU5noNUeqtL9m7MmOCZkcheboEEi+wF9HzQlCrhYPg8b6u
SgKqiQgm+GQ4fuOlZKQqRjZ4ScTEL7akJRXzW7Y5JGsneVuxV69ptJREiPmV2lzxaCJvr1GSqZ1D
tAdQTHyZsGjB8ZFD7ZW6eUPhLDWNsV8K/33Pe4TtSiuhLkrutU7e4XjN1I6q+0pF3TvcAayzBsOL
H1UPZ0PSlq1VELXnrPkZZ7UXEzayG0QT7Y338zsBplsSkdvVI+4S+tKma4YZ/OjLXtHeybQgV5N8
bHvZfZ3vFokHrE7r17vdhuZ3dh67BH9HfQZGQmUfX+1Bukt7AgcaETQpWD+ePjlTZwMBU3PH76KQ
3dpEM5HnDLU7T7UnZqI2hbxHMOAT0T0z4wxPtouWfzEAIrSDL6NYeXwBHTlT+3b1eRZA0xnuYfzN
tBxsGLmcAsELn7S02Min0jsWDoxcjfeZOzRxdC6vs4cUt2qSiXKTqzN3ydRAi+BHGrD0JHCFcyWx
Xej0biHjpLLL624/ePw8mV+PPHT3hXX4xOYbhqQgqcX26di1/UESBhHTEviPnZq8X52gWVgKsCyk
JZqL7iwqhKE7TR8Sw+B75vM/02KeE9VPprlbfTYd7pNdaPsFNHJf2wnNHa3JqYA+nweyTcRbrNGt
mvHfY5xBr83jwmTPq+qTsBosAuqkyMzIfXBIt5y+WG0w+O+sEcQp+ttiPT1Ko806gdVxLCllLlt0
OA+RBkea+4toIGOriLhr3IQzCZ2tEqyUa7doElUXTfo8c7sbs0SN7ycrs7FIFTHTUMWpLEZDZQH8
tk0hC8a55NlZBedpFXHYPeTafi/kgxCREqBmqJ/hoEObzP2TB0t55iEVJrmhUg89OgfCWLXgUmeX
thgSUkK/L/DeasuwGujv9hYuXFx7rc+DdKIfSbwxNS0qK3a/nvmtpodn8ZnAdK66CNDOjv4Wd2sh
ac0m5ID8VROSCDfN0EQqmc9NfojlB+Lm5aMgBkvZMPIRt+BD3/KK0iHvVkZ3gKPBoBitumwnLwFd
b5cbdup2QRNI6q803w5kuZRzSeuiqwF6aQNwVl1yb8Hrr1QKtHYv+C/h9JwRbsWaJZutmg6PZSys
JNePXf7ep9HRJRe5dThuHkz2yTxVckpUUMmjKK7vdeVWdQWS+qxs4RG4D7V8xG7RH8iHc5zYBMKm
NRrG+zfD4jzeOIxvqRNjR1KZm379dayFsJzz0dKInuDZkpDDH9fGhQ75gzy6fzo5w4mMQAs90rLT
hBW2OcVGE/ac7Z5ooqXHKgRY+zVwyENRd/zqzKLLPBBwzobS3G5Isp0oJTisdDAGpiX0D0oSXSiG
1IO1uGWnqwBP1q8F8Ypz55FGVdMNcHvngAqnOiPOsVRkC4kjntgIn/zRzvkaH/tyAiNPlQrTzFHo
apMdO/5nCUkf9R95nvtiZ5pKM4f6N3MIJrKaTOKDJfA6wniOnxUbRbhMt/sxaehvxSmmr1Gz42VZ
eiyPuLj/3Fug8at5pQWx7JnbxFOh30GMcau12GsDGj/UL+/vsVAzK/TZNtuoBKCdX7NtX4RMY25l
+BAbhrpnNe8WPVwOf11eVhehPa1SreIgaWOKcxWAAUp444zr1tCd6YGiqE8LVyAZOj+gDccRxRSf
Yyg2mZZZ4YW582F8APOF80BLNEiJYJ7MMT/WmkrBXopNEyL9EW++0pn3gvmdcWgPsRUi6ka9PM+n
vC18AmQZeD63us10ujf0xuAVAVm1PQXYHt/mJ/MBfCWvwvFBcElYvUAjCXG7Hcs7WxcyQxDebex/
xmVyfBUoc5Dh1Hzw0yUPzFzHFwZ46WbP1xwfHdv8rHgLzSbhBYl4BSh6L9bUTP1QJAgr17a/jMNJ
Lm4I6jKSTBeQRAIs5dksMgLHacqxW8HS+74fvYM4kA2bdFFlGz18sKlQhAQbs4pAG7UmWI10rxd2
hfD3A8Alxwnm6IDPeBX40xAJViGkUZ5+rR7k0xOT94dNYrkpK0k/ULm4OeGFWmsB4/F/AZ1OCIeN
EobCSoOTIJMRPcKsZzS5IB/0YA788pNu+MWmWGIYha/FLgrCrm3O8AZHTW9q0lYUxenmTnCTVUir
TVv7kRMcNzX6IWI7U52hLQlBm2MMkxLxfV8bjJrGyebYj//LHkpAK7VqoskU7nw6gLYrCywTmmGt
Qjb127qioT8vDKyBkPD6dYrA9Kelaf1Db8+w4N494MsRHusp5wlW+ftbFPPQ/HUW1vDAAsVS4+J/
GjYFilfVZJtfpSe8h1jERZ1eHrjVatBZhQJDuiPEn2O53MreDSGyXKKNZUEIwEkX4GRTtGTWXpip
AuWLfi39ULWoTwaM8/mneMSA2ny3DsSdPfD72i0lyunRPUDTgm4BCJvNcCxImqisNZd6t7O6hKdV
sXJRmSg7QEM25AuRAy4giHlMlGtLUEenSiXFr4r65Z6Er4k66GbZvLTd/H8VIcMQEQoIyXzP9ObC
ER9n+oaiHVnMshV7Li7RqHjw9OjyGronXjKlfshkKtR1yIf8Hfi9ODfk+Ok60FvTvG9zai+sSuvU
ewSXraON2mPtD3YgDVH73rB8xiRIPt/CFx/ocBbG5KvFfIr189l8pnLmvKqVf699fbK+5lAA2+JG
gzA9CT3OJgQeNtAmTIOvYawwJjQGZ9vP//statUraJOWcntF3un+wFcr3I3fDAQ8KoI8LyT+bO3m
Z8sfyKwDpRcDE0l9N030I6DX4tScyTYC2uUL1FxQixbCTbc5L+xHfoI5IAszz5BuWhjchCggekxQ
o7yI/a3NqFD1nzNZ1lvz9Qx6PC8beokAoEbP3+rnDFuoBhnyO5YjTYBTzZvzOixCoJ5lbfMIOrow
IMtgR/c3XwYApAZMVV0kLEWYOJQEYyOk8Jwh/NCs3hLbiuRFV6M+Q4cR9reM/e27myZyCQqW4kUV
GoQuNLXnkOUlqbEIJYszRJoYSdEYsh2YRzrYyvuCvXMiXxQf4Gz4WNo6RkJL9wESPt0lJGmUTDjs
F3HbzSD6a4R4Zt+tAhUVpJ2hAvrFbHMKDZwimtM0nv6WuaXU1SiGLYtb/Rq7E5NT99KhaNkyxw57
3L9ffU1gccnJyNqwlAKcFfAfV4BVl+vQaZbuDAYsirZBp+SSZ1Isvy8scbN5znKsbMw8kTVuLVCG
VkmxN/C1EUwrP9MwfZhroNu6tSI0jqI7jldbBM7x/4Dhb7QIt6UZPaE8iR/enp+X5AbnXt8Gaj1v
UVReA+mUNO21TycOWWWx9pU3IGhBYyhnmF6HsW7bjj3KYyBvLwbY04AOQ0fQ8JToiXmJfHzIWJxH
wth4sPAVi3JVzK+AXQ3+/6bbnBLOZdS2npX6JsmXrlopGp9rJMYgcc8QKQLg+A0FGu+ZKqOFkl5L
m2bj+6cgkg8UMcGTM2RkuSQSNuCKaF6NUiV9gCGM2S9snj0LdNLCTGaCVY2JozlurCP7ZQOd2SAy
sXTZ31ryOk5qHO9OX4500oSMYSRoQIn1fTAWNZsTiR4JAalqPqu8ABecKajjyf7QGKkm0vbuLntr
eTljY042VCTNLjPOvUfZqds8Zd/NJ58TK8xkkhiy3QPYTh4rABG2yy+XjM+lWhQGp8ZnDGgC3P/N
RmLtmD7uZF83kau1UjHQsA8RaS5QFUb7mF7feyMK7RcVOLvNLxDSgWSxobhF2sI6jPA1txpAIA6a
cU2jezU8FXtJAG0b3LcPZWsiJwnLlOIomViiHyO8vdJBAiuQ4OgdSMKC4WECVayR0RE9F3PBDj8R
r456PKXm95j4gGZXVHbOUJ968MOdG+YJbrVwkOhCdN0iO9BRq0uP8Bwt3KlAojEAqbHzxMkt2p9c
LFk42PgPYRBxOzV0ojcVuF8bSmnDFiv1IOoOQIn+Wb6IwBpE9P8yMATW00EydBftn+L0HXOyebod
OTMhRsvmdxOnXD/4IbgRyanaww+KMoGW1QcxXYvrWL9gxoMe3CrcDG3Uw3NI174aKMTdfXzatjTV
6LsEuQeDOEphymEUvI3GyJwZ/MHB6TwFvJ30TmbQ0TSXDp4lRRoDomwZdBtLMpGw5ch8MUmYESln
ZKTEZoNrnZDRtHg9QTk+40q0n+50bTeM9UP8KPhmo57vr2cAbajyh5tGjN+QfGqqcJx8ihje9b+e
JZJF6KGpH8n94JXx9Fx03051wntNLGyf+lxIiSgT6oSykv1v7ZTxGJQxO9vlP3MZroccVIrnv5/e
DPf+4A4djiZNVeiUkiEStRqImlSuwmDKJgQs7In7tnk+rUBJerODR+DJIwmF4rgwxNN+TC1n9zmc
BxXuZIu9swp85pwGhSLxwe/IX8n1Trc4SYVyJr64DKCNdiuurgx1KPq3kzJ5Bkyg6rjerLBvERmN
vt35WozyWkALXlzMbKDSCK9yHftqpEgCHBdWsaITJhOvf8MX2bIFU1xLe1cBH9Es0A+CbJo2eWSC
WmY9+Pwgo0aeNUnRTiBsm/Cs1d9zFNZ2A+P9Fktnkf282CdpGPytUZWFwfW33zlIl3BhKIMH+5+N
gXbm1NBL5nT9pdKkePZ1Ydu04m3MkAzJ8DW2JQ7gwwJBGHGpCpu9AoUWKVVWIm7rV/fPaPIMdafV
yzJaFIwD6c0Ga5acDpSlzMMGhPKIUZRJmqHNa8OJEFHmS3pQsm06qaTiunxJW2nY4d9RYkyKLtqm
YgmHsIsJOImp/rbYwCrBCSPJe8wHk77l1MfhST7PJ9eCHucNjt/Gl4h4p+ARnSgWOhBbgHT1NIqR
htSUsIa6m6OeM9HPlbdKjGDO4/3VbiJfqgJee4dvICLmAGbjXyaPcoGlYBxoS93lqvokqedy/xXQ
kwOJs0tehprXFkbibStanB5xnWTiqDShSdSf8qUrt4d+FTsV0ppm0N/7QH0q23iLG9w01mH7Ti+F
3NN0RZg14A6loLb/tRcVYQ7koUm14SzHoGqSdBLYDF4zNn6cm4MssadNckhBjS2KYQ5INw6dS2bO
EvfgcdAwReL+Y7K+4NI5NHpt0LxQr4Zgu3pfvLc+6PGai3imG/bnhSCIqDEcgtU+W4ks21hToML4
htMKmfpq+D8h//OPB1mdzTpmErmKHEM7ZtMjzSXcDzNBjGqiNJ+xEBUf7/JM44eXTW141uqKu9Ir
2F9H914NEw1jeuz6TeGSeHm2GT+iyhfazUAgvIFniOykMbvO2LyBeL1ejwwavTKoblSo7e9CW72z
+HO7oB418RuR/Q3wJVY7SwEth+aDj80nw0vEofT1CFnEiPrvAvsvizb8jRc286qL9rvja29ccUUo
9jTmCGqQ4grGyicxJMJij0tJPuTpHW6tfiuUh+fOQ5N3lQ58mJRZCFjmgbljiai9nWruqMO+LrrT
5RWZaPAbsp0760AZ9A+oXi0RirePRLWQbwK4qt472k0uIQ30iVCWJuZ3FMwtp2AsMcnrvubGRsFK
gfMY70eSmrNCDgJHKL+B9XbOjC4YI3+ssfpGQ0Wp1ZWmyQArIZYrosO5bJ6w8Lyvwqxxyo+KawPd
FZRhD2w1WjZ/1BU/6hYRtec0oeHRx+yBRtYfIjQfxGC46r3h5Dm8Ay+x9M9kbIh+8ye1sw+U2YNF
ribelJuCqhf31RDKyl9XLXAvbHf3WUesYNklFek3qN6NBKczSxdrg5Nw+kXlWVEUmSfYTuSZMQdV
OFc8LVT9L3gY0/LuSNkJ+cr3kBHgrZIf1Ft1APW/zqY0+9ESkuijEqGtbncswhMvxogRICjtmY5b
UeWBUdV7z4jeCf+/zOr1ZL79pZiigOdNxg8xB6Jryzu4jXDhh6n5mqDfn1WN+R+h3M21/uYiMZLM
11YfuREH18o6V3zMH3DWalFqLfUjvJCTxEprhSO4ENm4Krs9Qk+6Mh2h6pZCvtFg+XdVTWs3tcnv
+YY0EwhkNnjdlD273w/gNHxRsDrRU3D0AWHgkkEKdHrp0fIZSTJw3NXyQIF64z6DFevVazTVIxul
CXoRtdfcAUTwZCRGPnmhZEknn/9d4XkwDkDQjUABoOIamr2TgtTIhdA0qK2R1Nf8Zc1DNjAjgmVm
KooRWO1Y+wSakOSJqBFqgyhaZgypZaSTmClVk4Ku6HIOfWVGbJZGrLAlBuviJXwaYxNH493ve5OZ
bUVJtonAcpP9+Pg7TIGVCZ6uzs51bFvZWQtBk+Prco1I54Uht6ZjP9Yt8Wba/UlpT+/L/UXY5z3e
DDw4Ug92l2bkODXf/OxL9h8ENqwUXo1Ag4naxP002e150hdcAyXfXtRuL/l6XG0esA7mZ9Th7x/5
+7b0lvucWHsw4fGv4XbPLtvR3NIDNqRl9ImNL4yHHQTz2vAwJkg0c9xHmfLdH/BI5tbL6GpmQKzJ
xPrEzx3OVFjjVoCCE/cileP8ajIit1TWOnfOyFdKFrPxMktoUoF7g1VgzHhoXPBQT0z78tKUgZyT
csyCVYwAxEmAU+1lnajftG3KZeoMeMxw25p+btcxvIlK/p+fbBfqk+1b2WkUDaX5hBwqNryoMjln
2psqinzNBpGRb9E7kCPGe+iSXYBtFu+DmNTmt5lfRpuctZMUItEEGu/pOuxXDMW/4s01TdkgmU/B
kU44Wf3aW0j+rNhj7On4D0tjrRXYjCQFY5KjKDZNobpxTO7gg11MnDSC6tXy8TE9qgEfAuw+A5Fc
U5kTG43YZEn3LQ9PMfN6K0atw7oGiwEvvv/x+NdgZ9g9XMSfKpaZUTWKyJLaln+Z1wHVYzH5+Y1m
ttS0N5Wz+pLbAvGmTGugu10w969rpfxcFg6KWzs2Z91o1HnUg/gzML+gY+DnyOvPz+dLlx5NOI2/
5xlgUbK4HChV3znvpwk+OfkRf63xZ+kMIkaSnyvFOAq7Qek/8SOJYo5ZJkyEFaXIVdpv585HDeU4
M8kppwnT0a3ixz43M9R+IgNsbbMyKUPvGN+PYArxnUXUa4cILBdyFR5DTwBPBr/K2r9TCCqB9K74
/uZ35OTcccTLbb/THHYvzL9r99QMS753hWFDjLXuh/f6f8139lyPP+RsmRHuGAVun0ccP/WNLCW2
t49v03lq3cVy5ClzydVdqlcUnSdw2pS+UURcPC8h18gjigeoXFmvh99Eo7P5qezIsMs4C7zwy6Qm
6j7E0YAoALijynRiNabUOSGHrSCSMPJxxM+iDGDxTLO2+Bc6Py+es6MJgOofcowan4vo3XeJyGVw
e4dZq32i+h3bHfhKzFgGFHmPGUC4ljG31B606Soh5IOkpirn9XoZws/356OToSkh/vPbtkeUrZdd
mJaeKr/LeJ1YyGd0SeelHaI9F8pw7aVHf465OWvV87nSt3uGmTc4ktdxNGZXvYPyTpjg27m3pkjj
ObEk/1nw05mTmihhzJXLye957NyNw6GB2Vg+m1b8GBCNBQ+75btS2eOQNKzuwp7vFTxUhn1GE/yD
5nYVCSqk66skZRocLPhaWAYhcfzcrWcmj3W9UkYK99wz0JYI4pk372nHYvM2pZPWmy5CqCiSyDZ3
oskNZR+s+vkqugYNw1ioz58HAWIU10gMZgupoUWyqpawwvqiTwDZ2pqiZWqTRYJe5U3VROLjpZFW
KS+1468jF1Hcr/3NswrJvsvQhFb3+nqxpMOd8tu6eD9qOLE8G+YTUXuPX+V0alKmQwcifoww/k4C
HyR6lFD6Fhp4jJ+0OUG2/cVknRKFz5Kt9Gcxs9H7yhHPIgp98i5uF1TMZ2zFggGt/lawGqw9GJ9K
T3rFUXUPGd2pI8fi3zgeRArasoBQo1yF6GPIlZ/MgYKh+rEUA7EGzmKtqxMrtjaQED22JLkVRvly
d2Z72MjrkUurZvOIIGQxwFjT1ExLpZTgH0I+QxCnon52nUDMt2u4w0rRBuVGUQOPuF4CZDs5BmWz
2jzqbYzb4KPP1UfVAp3CxkEb2CxVMgIxyr0G2hwlaHBaj3FeVs6GVNyJQR3L9uCgKzHY7JEpcs6X
N8noj6fZV7RCuL9NYMe8ShTGMicLkX3ZMe+WgAsvdw443oVMKX4eU0HXX09iky/5X+AwW2cEWPiR
zknYtHtdZOF2PCZI5/aF/QOCE5av70MQm7E6F2q8GXK5HnV0fBX7AyJK4u3iPUb8qa0OkTKsm2Td
EFrvuHSKtXM/+eB1QLcRtgCcDs8aDp5AtLVPnFMPvYUr9armjdK20hxmKbDWqCWIPkjhX8qt0UHM
wDr9LoJU96LoqxaQuKOdRtlumV8krfGnJODaJMWVpvEm5r3OcZZlAO54s27f26sPfdgHGWVx4h9Q
h0mux8W+FrIFcjgWgH62ne3PDfbVrT1OfOXWoRBZ/JgyKXoGapZXahS+8etoHz3Rh7o/4QKgN++Q
i9EV1pPvJZXQ9e8dnY2TjT8Q5z7DOMrMUOmXarhPxSpffkYT6+Ds0wkwivcqjZdrS6MrshlXFcWi
t5kN1U1eb9Hw9jEr7t4rXAIdnfJ72mxPaUoIfVMQf771txTX7nSjuRFoM5jOS/vDcXGKN6dPwHdj
G75mB7j0zMZbk1NIUBohHewT7hW0uadbCAKOZH6jbwBHoBAkdymlWrOhOvIKtoh8Eh8GN+JrNQOO
15EMQc3/PhuS9siKVL5QjDdd8zC9E++J9m7Na2YaU33scpZJefVLlBd2/Z9XNd06YBoRkSxRpnXf
iLTEI6TxiFbY66k5Q5yLU1BQg5A99/1q9z7QJvoK/VzjJx290eMG+aXs9RL808uy5s1qBH/jtHJ1
HM6iPOZgpx0XYp6MsdsbKD+YZAXJIKSdew3QN9h6Z6pPA5kcemYMCwpkvI9lfFluL6BbpirwW8uT
jwAgy+uazshQpsuu2C3Tf8+ZDpxy+/p8dCDNz5O7pZ+fDHyMF758wfQXnhZswQQjij9dfV3IIc7y
NTgsqTpaMF+H9GTyJRcns3zl7kXCivUUhoq0XuHFUUCKjZH7LUW6xBTwtawsMcMtzfaKOv0exD+i
Ik6lKlThyfUBF0+os5pLjTDfzGOAdBo1u251aN4OT4xrWNqiQ47jkgm9dDAasSsoNtnMV2uoqkQm
GSSSbeNANow83vLxnrEiAHC+YYrRaAnnP/vXNpVUaQsPaxrGgLFI5WORgNVvrd3TmCaym5GMp2zz
NNl6i+6S4W/3kzHS26FhMWa4hMm0mUiaBiwsZD4pgMsC0hco2wYRBm3fk5h9ePf3tUAfIMHy+NgC
pDHobVdX2c4maFWkuKqnezCGVS/bACESIm95EQEmto9zeWyzT9XTcSZZGuzk1VoYoJW6XJmLD/NW
GjkLfxLEWDrG2C+bSJFFOQ5675cD8yx2Xu5MaC2rQEdL3nNp1e5+bC55HRt7wjWhuVnTVGf9keCv
Tm6u3MWFnFOu5s8FIxoeoXT/7KFPMlz0CG9c8S1ClZGAtI0292lkkJm4xJYP+2JqGhLpmP9X3A2Z
Jxox3traAeZ8drFOIUlg0UpVXOkaRAc9F1j1QjPnhD1peNcqwC5v/eaGQEyPrfKOb84ttszCPZKU
w5QNRe6dF69aUoROLWG4AE/aQ4tkOh3WkoX8CaHNosTmA+ByFqATbwTyI1lT2wyHWS3a0oRlCrRm
DbS9EOLYikwGjjYCe9Ujbce8dmR0rNMY2k8uTOusXOSrLbJ7cMsiyPTpUF4by3g9j0dC+Af+qRce
qYv7XjpSAr0G4riSnfc7aSgzEYoSyCLIk7uXlNdpRMk3i5VKkuauWkgN/B96KGz7J8jX8oabB3px
qv+lA0qceUXbfqv2u7zVLTaTnNX4MCXRUyvyhB10BjVeCACftlMG+GZygeYWSo+KfnbGiqfNt56j
2wagnloeeIaRh/eDURdrnsWkYkFkLIxxVbiYrmr8GMhrDysMuWEjxlFpo1p7FabTJV8VtiA5VRVv
FJj9itSPUYtkQx6P2xEBgei/fLtjs/btgGf9Vq2FE7i1Y/QDjdpJFPyZSWPBHr+yPsoZCuvin6kA
m2vqEDJjdQbzl3eNVuV2bCx3/Y7dWD3gp5sUl360HJEpSJbdKwdwT1UTGQaa8v4SYP+IZJRiXGrM
vhebFXcMFPzoOi5qF0V57+TNIxHyJ5Cackac+mu9rENgDUYNtpC2JRxuKEj9Okq3xLvvAxuUPTzn
D2vS/SakdKBlcFifF5j1WulK4EAVeXcLXNcv61QVQzSauIJ07yWe0awuLt7MSraY2oMGz/B/2WDd
ljPeskGtbk9A0Uu64H/xngFaqY5H9f33/yoUsVOY2wUMfrJ4WIulkT5LEhmit0AhwDSmDZAW/w71
mU4M7G0UrWrY8oz/U7ATzyO7559xynzUEzY0RvVu78vvvame09v4usiANZtn35i1Ei4lI76zrPo0
PvCM4IN76DC+sITzqrB6tL8+Ep7EnbTn48Yv9J2zIG+Nzpk+fc7CADeJq5icK+5cv0LePBXT3qXx
eAk97RoOZoFr76lhYgCs6EUL6L89/JyafzZB00GLX+tkCI1iPV8SzC/ueO+OKja/LiuAp/3pFdC7
L7+eaAObRq2UoRaXL1ry36cJ5a/38sAtiio4+JXYVd9mRrIz53w1SEEJjJqn6vFjUWE65qcjfYhP
u2gjODnZO/1sgfiN3hHE4go2H8zCf/Zqr6UZy3KdKym1dqRcoq0WcjzZavxlicRERRLCzRSzNVbs
9QcDILNhYke5V9JZesnAzdp/QewFXuYF9BuCL7PEDZ/YqDbJA/Kw6IqbYCuD5s+C9k9Ao2Vz2JNS
Ni0zy9s4zZGxrkQ92ZlQSB8zCfEtS1FNG/6VN6rAAS+dwFwov5pxsKvDg46VWVID1UHR1V0OfBOt
HExFNfTEs3Pm+/f0Jmj1feqBPbBmJJ79Gv2+d201wG/c2vLdkZ4icq5SLg7zAIz9zmJUtgOoSXf2
uKINcljjEDePSml77VTQ1q7mr392JF3SQNh5SGFsusM5ICcE0upH9gNrzLZ0+hl/xN6Y67/ACBSJ
vW5z/1ufnb/5HcT3vx5b9TfoiatwbbT3oDt5kW0pws7LZcyRU2KTgzfjzOV9mnisvpsJBoSYkW7r
sHswpNgrvDYk/+q71T8Gd+b/72vlJPMfZ4j/Ufi114mz7zEnpqrYx18ywd2vSXjq0cdJD/FCbO0F
KX6JuPkbETgBAuqIasDYrDIASCYArP4Wy38hgwYdW70FmtEWQhmoVX/h5vgIvZwwI/D0Ad2I74Ec
XFtAa37ZnxWYjytDERWKQh/xOzCZflRwBJ8qZe487SIDrB6IdUyrnlNqRlrBRpnbImqn/dpZ5FHx
9fJ7pmzLafFW/84nemiPwjCCKNEXadXRCuam09aLVYinBCMfIOMFjXM/YwoClIEwTxdZAG35Rofl
alU/GNm0d9GN+eA5NwBL/aBn+r7W1fqsH2SgerYDzU0mTiwuuKIb1ijXSVFRidtpQ48CMwr3ThSR
EMwPAlUx8q7nvAwD/+33HtEzK7teYZO9cMg8TbhF+FHBIJLNjJoA2nndbhmzliVM/7shrHB0dfQ8
fcBY4fsJRRj46YHB0+RGnhlTVc8fdFytGggPZgFf+R9M3DPx/3g3yH68pnTa2MjT6KorZQ1C9jCp
NvrU0bYXojQYMp5OshLelB7eATyU9HYNuuyunFfCxraUx7N2ljIyfI2GdtWakczqJGOiRvPRfNea
AmueyXXWOYLiSbw5bEDwf/AYu4u60HEdE2kujiHGdNJSg7tTLgksteCHwjyO3pAGaMoCHyg93zUL
mKI1gMTih8JC1k9v6APdbl4NLVGru8wchR8fo4t9PkTKGt1g7h8W+Ll48edTZ7aQTZWl+rOc8+qP
5yaHCqV9aUAyt0b525gbwVDGeJjBmJ46LMHvzN97m3/B/+0kCxoAOlcRaj+yfr5UOCAM3vz8n/q9
RBWks3m8P28PcHioRUb5wArgCH7sLMxcZoXMkATrBiz2knvCtT9HlStxVnR7xxV9rQ1IS5unWuJm
QF0t8S11DHCRZtajaPcDbDnhnlcwTa2EUTCspUMlu029QGZbhKu5/er3QqnwHkeKz896skUPoMCI
R8Gma4Gri5pJ9gMvdMkhP6EVUhqynM37JKv6HcOLrB1FNCxJFIjDbaYHBS0Kt5sPg+lBHn+fYth7
dzCyDwT38LnCGGHYEMBg5gF8kqUsavbI/gx8HKuJoaCyiXRtmN9TAKuPab9CY58TByT4D8flTgzi
jhphwSVKwcCO35R7IUeYhbpLYHbmC8hzyo0wfGnA5ve/44uKOr1Q5JVa/xlqeFsxmIqkhDwWAaO4
RriDl0X9WCBcQGO/aHChecn8U9Oer1hSZM4SLsBxZzsvaV9DMWZ+1A5WvNCtWFKfqXa4JtkHh9tk
qOo4ywCbZNrNfucqAyvos1YwDgEY43wWUqMY1/yNXbHs8H6SmFh800rfqm9gdLFRwm5NYmBxHGBk
jGVqVJ2UIAHHaZ2Q9j4gLvO+MoJIXzRyxARZz4hSvbgHPObUcJEdwTBEUdnDghDb+F5xDB/RspA3
ep+lMh1Gj91s9t5NpbEmnDZvIqPINTfCOJgkOxoLKI1RpJw6yLR1DbJBWKQgrxE15hK/rqoWqrXg
HuXKq+pTkbtgb8O4WivRH9F4cMfHvqG5gD15tRs235Qr6kpWggyF8M9Cf0zajj+9bYWVdK2YXfCQ
FXNN7A+BpFBDDkS/MPF2Ae34ZrnZ4Fcf955HKHJKowx5C9fb87lVIY/G3cxvR526GbSdJnZj61Xe
5y1WjihPKaC60TEbzTEnhf1JaIPMi57sl+BSN6qaOXe4J+DFRQtWAb3LX2spqcJT2SamyrzumLTt
hCjqYFycmB0hglrUOfLeEBSw5E/hrJFByhfQR0xvNN/++BGu8rVoxQAVIkztXr34/q7DJ1G8MroQ
vs4WaL7wy5l0wtGRRBzooyoA9lDy2kBxwMijjYuFzBB54fnoNJ8hAZ6S0iTvOegUzXL0Qn+h9nTY
uF2dxBSPcF5d0xFLIMKQuX93faAJ33JpZUDXhn+4F21QcxRxZEW3ubUNj8tL2fO02ax8JFEzS4Hq
7Sg25M+Qwt2fixuLg5+gjBoThEYOYrxsRli07TuMQhFA5ZSQpncNTDbwfAsPgGRcVBKKoKHJmJgM
xP0p+GDrT+iskY6tMvTBf+0mX0R+hQ7vldjBFJkSBvygtnnwNi3G+FHYqtjfAVCeCIOUjbz/HdyE
Nl6XAyIY/ZLnTGUy8Dm6ZtCB3wKKVPR1WkC7+naCu80FhI0wi3vagew7XvM/O3BP6gRqsHZjArCP
Q67Pif2cAelxeapgUXvXt4xAWiQvrG36ANZupo/2ZGw0yJYPexJz/AnU2FtJIthcmKxwGD5AUewL
acAgvDFgpnehlCuGrI7l5YMNVYODwmNUvAX5kWw69jpT5NmKzqKgT4hmNJNtiMfxILRby62wlkDv
3X5jFpVZPc5wmUvHz3rAtr+LR2z+61SGdniswb9OtH7j7T/4EamgAIHt2SOKUV3rbcH4elXSQHf3
E/PLM181lh9ttouVwS7c/4ltsgOiuXq++8L+9E4JS0opo0XYu4KZpcQrqbEb1cDmg1vI+9zhKtM9
OG7O0dea5KhY+fvCMaYoCi9w/KT4U53s3PN/ggkcHXXJ3ueFcSyuOVFKrCDzvZ6mHVfATDGiBlNf
4jOcnJu6fX5HJhEGn0uBS+LABEnakTOKnwHSZidp9+VsFGzctfNBFu+dx7F5MPPgVk+LX0IFg/TC
w5+JWpTb9z/wsXTSStDoTgEOAL7AHqjlM2Hy53QIaDHi/L4ft1qHkutR7+VjKMNqms1iR9i3gXCU
UUxxF4kXRv+c/eZskR2fly7SX1ZBGab8LRLdPstUn0OEpDu7yJS79jUQO3t3J6EcWQrizDaVwgBE
TlejJsvF5oWbfzL2//O8/hBGZpE0VvqrrL+iLeikyyRIgnQS6GOnm7m5xNMHlqXalvOzS1SFM64z
G9HcOmu+vlzPvWcct0hS3MRa7E3Zscj4vvD+JA5dFE6XNFZTof93p/lAd/ii5hCYDp2xfguewIee
5uVEeqOUKNAcO/b867DVT1k72k1VVenX6zSvB5rY2ikzG7ARfiV4jC0/ArQCV8SUGYGL0lzlBnN7
OijO7Ihiw71DbWRjhXJbc+5OGNJGdWCEGI8zCQJOEiAc4ygMGA2ViNIjdz2zUvnISgGc/9k89TuT
9QB1BO/u2s8p5uKBcqv6mZ84LuDzgPZLA8+MLYxQVBTHKzRy36BbuUC2iCfq2mmkU3aptovuvQ4H
BlX1u8TeTfukqFI6XB3gWtUDYVxqeH0msmq8MaUzx67b3O1KkdSIPPjDLz2cEtPPKWAnX6kOtUKN
9Goa7+N5/z/x3Xsbo8346aSGF8XjVaPD7sqgTuUOEuur3cxFEMZD5mx2sYQz0TqZy4jbqtVB6pmL
B18BewU/m/YtueAX9Brlo2hEhxqt4bXMBTO7Wp/asuUqU77pfXfXgPkIbLRv3xHlrEPvJsg4PjXR
o+baAN9tJxqFE9F5rpyYvPJ4jSr/VmfpT/ZnFKhV7q957uh8eDG7aEN656fT641Psp4ZC3Te/1QK
fyGFKJG33euCAwwO0SN3SAU2agxkVwEZzKmE7qTTYXZQPJrqFkMc3QWzjaLDTuahyFcNHbPrb2vI
13kSwDqhM5ne6qzb6Nym2owu+lgyOxn8NnnOK391TEWptCjcolSe5DHslE4Z4euey5K/A4KJYpbA
rxRKSlakFV2bHmzfBwQEMqJA709aMiRVFkLFkKgMMiXtuFPRctU9dRWJxGPt23y3yuU68YqKwsNh
+wiErXZGZVG4GXDY/ZgSTD38KcVlS8204a6OuXQF4vfR2fuuL+Y63sdpvi+Gti/zF43AWibzsWmL
daT9WeU+FVJ4bh1dEh6+1B9LpzFX/5fVjNqQgXt774IfDvBl7if8sGHjtFIoEixzPhGn9AQLdW0N
Qc4R7fKYGCFKnTuE7jJ/Qf3pofg/f1xNP2XfreDZawf33kCup7U+FdZ7bNsGStDFlV11q5MghzCk
e2LI+dml5dzSEkiWhZikyxrbAaB5Am8R0ENpcAHczkrF7f5/3X5iKAvmiqUAiwpZEBC0waFaYIn0
MvCx5GgVWmw/xZWOcCYu2FNDmCZ7PfLCKRQMhQQ8ZWBF1gBjpil69nwyWtwUekIMPnxv4LjNP0RC
mkfeoKe/j7ZruS3gulQW797mmz3rqGBEP8er4Uj1SYBk+Y7aA3FHdJRwh9qxQVira3ObFrxQwTC0
PJmPx4UxasgDVapLfuncdAQX5mSj+mFXhjLta6J/pzDPARQp0BBAp16jjhfTQRkXf+D7/knmvRdy
V7GoJT89ZejdznvvwKEkJ7jaF+qa0p0sU9tOgBpB5jDWxP+Jl5qF1sUBrHtWdAFA5a5pr9R18Zaa
j7IxZZkmpCwxjHYeKRlEnBUUHMpoNP+rqrqXaLynOFyePHw7Cx31GjmbEBXy3YchdKN2s/xwU5qq
PoZGZb5vKUZQArljb+LOliPN/83aZufpSWA/IBJSwG9xF49MbNmxliUUEGbdMb0arDlZ3R2IgFat
nwLaVRJjzS2ExbMBMpLWMSYVeQo/laiygWkmhG/NS3dRO/GVBxiOuuYFM/t8X6udTQRcaqyhWEfh
cqv5dQqGr7Qw7CIFH+XzH3BJbfdwTNQJXkIkoXSxIr1YCwIyiCV0DkuyfokSzBzdOAw7dO/zeO5z
QU4Gia5fJD05aOzA3QoZ0/JplUP35cW1+WiK9wGdKnaNiz6XOthqmsHYIgshpoxy1RaQsoyOw+oP
QqGtyak9uF4pzRUzzllECcQmi0iqy/VQpeZI8AD/FVon5gBf0Tz2qZMZVOO4+3vhQqfIg69SM3LE
aWDPeGR0HR393reeU17MXR2myRh6warvKIHLvWBaSPPSUfX0MC0verkj9IFEydzfsonSzlhMSfDx
eJCv/rYhd3BsjsN1cmOKbpzbcYT4XB4TbRAdMi2Vl3QN6gr/LP5T4AGbN+OE4wIg2iRVhy+Q5R2a
+Bv0Kw4+tOTqpqLemUVgV70vbsbOh/lr87kx/QB4UhQJGkUo4NkR0yc7Na+GrISZNqX6n+X4fCZk
xZ0JjwUvjq0pq4+2TJ1WZd2/Mq5MFHu5wbDcE/tsX/zBPhtXNrN2SGVb3t+/JurHhm5eQtWvWZ5k
Oh62Ly81fOQEAYujaJ0WWrsrmbleSPcrAaQJVk4UTFmRYsZZSkuf3Lb4uyO/4BawxtSYOsxa9J5A
3+EkeruM/6YCzxBhsRbkmf435LfHvuVszHlSL25FvifhzV3TJsBwXPwQCt+rJYxu9QHO+WsQPlt6
VPcbVfPLERjWQ0y1CwN+IjgjucI+ZCfiqnZq40BcxKUCK2GvCDmnMbKyUTq57pqfJB+n0rXrQYKG
p5Z65cS3Qxk+4L09LVX1qeytv8b6wBIuuN5CE56yFOjUkDpzUccpW/dv+0Xgw2DHUS9eN3wEoTUy
q2U6VW+gaJTwADgWLTPcfWCjyFpAzmerM/hcPBcX9xm33riLPs1uen2BKikpFjWByobYRYfKySlc
+m4x0N+ofASNYyKgqmC/+xFwJqdAE+vdomoF2ADRMT1CK6dj/yPZbosT/uvjFX8YGuYZ0T4jUAYw
s17mfUbSf+HZAZlsEH0HmpWSKkTCwQfN3f3+hkAWjTTYbcCl+A7vuWCn+3G/kG7xOH9oB7cekL4Q
k+UnJ1IENvZzn+xBynk5FFi+zSGtDksQkn7CqewCYrtLOzJN1jbE5xw/Anc7NEffkxMTc9f2UXio
AZckdX7yPvHDqpoJdMZAjFZT+BvVGn00r8iaBfVyL9UGUT2wrHg7SSRDjVZ2t78DFWM7Z5rKTqJ/
a9baPv2LRyOr4ER2A0RWGxNvihUUDWGYGUf9axYJQLxM6I70umt9pOk2B2XlN7hUizU87TEcHKXW
uDN0FLAUi+wW3FKdPwl770sRg01LYaZafvc9wy8kfn+nlQpx92B9E7GwY7F7QQUH8uKFlV+U1sDM
obgnqp3QCk0DNQjy8SCQeXXIPrxoNhHXDw/R7Zdl1QdQZChBDU0L49i5+eNq5jL2+HEj7fm5hKu9
Xr2NQjgZMSVLv6iCFNzJARZTjHX6i7G+jDuGovCsieP2TKlFX7Pl6oKYawjCD2HN9DXlagDo5aCU
3z2DCsgV6yMTvcPoiYIp4nmgZjBRdWzbAJtwhzSSQMai/clQmxwXw97XGD5Ek751KY87SFL5//D5
9OIs6zOff+TV6252m5yUMvN1kmwrFpuvTLeTBDHWi4itD7dUfqbPoSQ49pDpGB6qgmxNVPNCpedR
6fVeuTMON7LYj40zxUnkYC/P902w0qw33mkieS39Y/933AKD8f5K7anXL2y5lYtNvd5zVGQh/UzH
he8qpHl7JmE9Z5A/7lcJtk0wzsB4zu/qhTVBFYEZI6zraUw1eja/eVynAtgPnfkx/w29aLcMiIPO
rubOOFIgKssjurId5Asp68D7vNDDlWC7+NBhlwV3B4MH7wbzH5/BIR/34XbyQ1JoTS/AVy4jEVE3
u1zKX2mp39SGuR2avIgYdGZahm0fobz4cSNVzR55orp1j2fQ66UixWj/pyjNLDmHEwS+p11xoLCD
yWyMIn6AIcy7Yhzth8iomIzzjII0jv6e66WFqfcHNro50g/FRRpamRoCYlOMo8FIAFzHh74o5TjJ
qQ7CTyeeToVqNKPdV9B4yON67/pR0RtPMJ4zOZrR4/MwfcgH4TQbbSJOIHxpT7gARRoAqrk6KGbS
bkgdXVyerqXr8HAgJK/ldjAdYc3k4RfjGdYXZQ/ngGGLz0DyLbC5XDkA6LD392PQBjE/PVp3p3Fz
xXcLfhLUHK1TIdgoilZn0szuf0UgOYL6bPbi119Z3DDLpZe8ZwIIgPpnTOUx48ARo/k0nP0UsDIS
YZ7eVi6eLxgmNUC6eBK5w6mPJB0bp052VKl8B3XCDrWxJQc7pSn5GyBzTYPwea3QhL7D3XBtZBlV
gT63p8yTejLKs5T8Y/LL78ULDhvAKV02WpdrhqKgO1b25gPi3dN+TB7SO0kpKCmhdZFfXsJnIZ2B
cAh8mhHSDRMIUFx2W6Bo106wWccNfsEMY9pFvw9BkebjQqba1hlfTDA87Ck010gb6MSslqE3PUVg
5uxysLyDH1BVtB9ZFHt9MGdt0dcorpZ4m/KCtpiv1YDI5UsU858z27AE2O/wDlzGTFw1A/DfNfuB
VhFNoo//Ue+zftwJS38cfoBtahrMPoCY0kzFxIEOhUg5x071A+O3CJsJ87SPTQgqvE/Pn0CHC4e6
8/IGEPTagbLgjDnBfBes6Lr/EqUdlLM/Um6kRGfaTaqYngRXLdv4Ny7E2UGpQb7oRJtq0hTIWim1
cYrqzcxFIE3lFD5dMS1j40BH03NrUw0vAQWY+ws3Xs6+wCNgO53QcxTszZP6PmJzmSepdO1HEYTi
ukgF0g2+ILrij9D4K+Lu9dPii/QovtZBkKnCPf+tdbATsvQ1On7Aqph5StH6n2hynM2VCF7x4ua5
E2ehc85+da749V5SWGJQpclFvxaHEZzdjvylWEfkoUG6xACUBfioxmn+xZniNToMAUENQKULCE/n
+55VqOKBSRDEL6n08+IO6GNHabqjClQTVBDe52pEvc9+Se0YSwp6Hc8PxKpRAuc0bE+q5YuoI4x0
cwQImwSAgx0CKG8gb48dml0uUzbTvTO8sCVMztTpsDwpx7/EqtjNfQ4C4xQmRERlppm272oE4BVw
jT4v5aDp+mNljzImbL+bewR8eWijmDCq5pXfgyESfo+4QZfu5q5SUsvAatwc/6wXQvigsS/tGGew
sT7qYwoKV/Og8DPi65IqRQeyJWvyrFbZDW1qX97o3DHzKQsRPMEICITC5N1pcTzrP7annghXM2mF
bKaFpCy+I9i1sVkubwgQDWXLz3FOzbTUqtnv2lS82c3KIPMUUFXobUfvuCTx9clIKBCr45lai6bF
Zlr1kvJtSR70vLVj3H545kuC+Xyb3/oJfiXZF3l9O+tPfHezOWEcaic8ennbQi+wxk8OVNm5HS5g
Z14MvCajiX8ipn4Asxotv5RxFEE8OVMk/2XY670F4QPyaIvX1VjCN94iAL4E5Sc0t2bYmkOlXvyV
A2FoxpGgcRKxmTgmM1hb6IZTZyVbad2FC7QiHNV0RX2uzlUbESJUtULTqm3MVzgFdmzaKvst922R
uaxPo+zdaJPkcGoi/9qxJyKOqZUUetVSA6RqPIhZOku7CGuMmNelopb7UInGM3de/MCDFVwK3mIL
1Njb+PVUsHhs3WtcVuSU+59kChJ1OB6hggiFqvgrG13TUjVPgjpgS3waKcobKLtfZGgNdSTIa8EW
iLskwHccf4LaD3baMj6VBXa9yTu2+yu9nycO6+X7U1HDraJZ9X/NGRhYSx4yDfWt5uKVdL3PuHLn
mD+ZOYRvDLV2wml9yHkbyXfAVuX04svOke09h4v/Q2jxB/nGvcWKB5K54rZaLaV4TsThRWWq5+9v
sG39u1DSAbSRmwswkVXagUPvI3Y2j/PHorsw4RGbpMadw1BUwAKwhlz5tKxkY6FY+Yu1oDPeOu40
tcNnjrKIlR2fHLz9oZn8lgzqxVOvX7ik7SBBYrzBtybgnx2UGn1fcYDQa4AGBJNUj+qT4DBVPqyE
18iAMxCOJ46Zi8Umck9/WRCEEemRd09kmquW4VDyrSO8Jvy0ABrQDoRWfBNWActv/jA2fvQm5dn5
6dzpl0CDuZOXcpDD5maAC8kt3Q6HII890KnsIKCpN3OWMLKvGcqEY42wZnOLXWY5rkkU9Cw+8tBt
X4zzL5gr4FNUX+pWGG0mjD0aoi9hiqWmzTMuL8It0Zgplx7Jkiy/uMJe2E10lGl9AM0wdk62aAsE
TRqA+YBbOSNewBzSiuvd9PIocHXNvrHF3uCP+8gyAlxdTCZVpyONztiA6uvSD6kXoZGGjqGlGlpu
HpLcMCGuYyACXxhJQhpl1Zo+Pjd5YKRlbSw18MZ7OjC/3pwoeTsJmodbPAFMvwmMInFfcUtdY0s3
BGEegYS2kFrxjJ8ygauKfwe9+/MNrcdeWVGLIDe2i1scvo1kFz80QPSQ8egH4cSGilkaMdyT9N9U
fZYzPJKMdu+IPQ2REhWhcS6rZsOl26N6jfRKKACaM4fgf9gqQk+KrA3QWjrewtiTmpwwcwuhsSh9
rqp8GEe5gbReW6Cq9kszAZRRASMfZJRHjtqUJ2o4lrXGDAHflqC+elswK3MpEMagEXB18ixcj9pn
phcoPm1OIcStlQffvIhtJH4RV21rev9UL4zMs9CL4+VdbjKTEv0tEXHGHywhYyt0D7kTiG+cBnE7
GnbyMM2WAb+3TT6gu0Bwfk110Nge9PuEdbEwfuCaYV4XKawYWLf0G6eSJcXIsCsD+DBUiGjBFMSg
GdGBfBatxNbdn1/WEHwUysGltvk7DUbXl7NHBkCjLcR9lwvEUtBBQxOiCyVG+1phBpHIynvfi6b2
rHubGs517N/6cm/YOemzS/YUEXmLdgV6aOWJ7J9zEZsDufzpqL3KcV0em9py7xvPjbZLb7BUk6lP
u9xXrL03T36i4AFiEbyXm7xrQj7GySkjMU8qfm4gg0neYmvGjdTwn+etagJupjwEsNrJJJzY5Ogi
UFODqoPAVV6M1ecj6nPYOGwK0+E1iCQe89/m14/2Iyg1GEzw2mfn0RpEGF7qiKMPpHmU3Lu/VB9l
XmIn2FtXUUFN45xtUzvZ2Klr3gieeU2SqNCHGhBXRb+aVd3KaxyElogeAfJXkP6fIlfYg0IDc66R
8k0o3uWcnwQF0bw1glqHrar0AWMONhbmTzFPjD0hs6HZgMzY0+phK6pjggYptbRPAd2eK/xuFHaj
e5FDQOVXyGQxD14gF006ZVDa6xytHmFYpLFT71qvVIK2d6fj+JFyo/Z6bVcDgWdDHMKQ3ae4qBHw
F/51SLU6xKt+uWSV92/TGiH4aYKw4/Hq0sO8qn0HymbmR6IvoDfexw+3XpHsFMJsCH68jeT+M4Qa
JpgYNrCleVz0xPaS15DyljaYkcqXGEg4lJbeiLoKCeMpQSXjUWeKW5OICDNJiYZx4gO6BjMVjp/p
qxaEUMHc7If+mMmBRojz8RxGj7TGIuy0dWXFKTdEZxkzFiKSNOZevzUKJxFEvCB+MDGML4RXzqy8
c9zYFRmNvelbqP6rJbVUnW51fTYdgmIFBOMlY8TOujPo06tz2a65lS2Apdd3NJrk9kxLFKqo61GN
zUCVdnUC2W6TC+fAR/HwrAJmnV//6twpgRcTzuGsPJMtg4jLX1NdvT+jDjRShUx8K/TUKN3RBuv2
cvvoHsMh+AHIyKNij42H4yaZ2mu4dnTFCLBsJgBSkOeXt8id/mih2DGD7nkr97BGF7pH7mTv/Bnn
K70tAyDu4o06Pk1yHZUaq1AXaAihbm7onnpOswJGerK29jmOaLWYOIjksCPZ4cSXWrsw0lMLD6+/
uQAxnB/m7LHJ3/g5YtWcjKQBKAlsoGFX4krZj6dnuNQ6xBX0FJiTKDFWtkjHmwwc4nmA3dBkDqI5
2HjcO5+zo1fJZlob3KS/bM+XPbaaVf2cTKn4+8KAGw53T7H6CDmvw3pXHaQlcQnAmrUk96pxSAhj
5X7VotmgYauaO/p0U2X50BEkMYIpm/jzkpVnrYf7AtAd8piUcLGxEuY8sJnV6SODWmGZf7gO1/5v
g0zQLgOmxlhjoaVgGdKRXimr8OKYn6WRz/3i4KogBPkP3iNWxQf/TQnHBGqyetJgNYNE59KrrQHX
pN9RHDc9zfIKPb69rbJPvBeBbpD1apRFiZJfFPEr5elnf/2h6MuJ8RGK34LVVIyOOaGL4cn46ldo
EpbGsw4H/4LAxuxS3sahU+P88t+TPEuhtkZhngfiOlEiHwBk0lk3C9hhtjEx+tmaj+EKyNB2Uli9
7pykc/cQzyQa6ytxYvpkmjXT/KSDlWCG6xgAYBRxPdIyigz8fMwji54hqp3lpFG2S1Wc62LiEJoT
Y2m/udJAkOEi/vG969rQ07FyCUovrPI8Fy2TY9JUljWuBDprg20k9si9bC0dBJivtfBiIu1EP55V
5SZf7I1s15as9mu3UvTo08wLwzzyFBUaYy0Ic7wCzaG3M6mCAvx7xO4FDR7O8FsG8DQdQ6cvsL/s
pjwKwq6+q6Xk5iznJU39drj7+QJzFAr27w/ezBL+z+2ZrF5BI79eJmOTQQG9dCaHl9xQG3FXHDHi
ubxf+uzQKKgj/C0fNtXIk0XIdKImdABLqZAUQoSDgCfkFqglAL0/RugwUQaHL6dPB/JEub866axO
+FRwX7JRPysv3DC6nbQtMNwlPO4F+N8fxWonxIC3Lp8qzlt4EM2ez8q6VUCELTBz9Vbq+nEagaDt
Uyp3DOF5RiMK/2E5Vkhp75qmjUI4U1xAaIYOb69iDZuD+2bgtdmrXEYIZhn3muH1ZdnjSb43s/tS
/+RYM7qWSZR0DmiHGn4bweRsk5iWxThYfmC6zpl7F4bwGVCi7akfoFfqwTxj+Pg4T5kYJirqK36v
DyQeY+T+asEizpUMEs9v/K32ZvhtGrY0+8WQ71ygX1/YkY68W4NDvXFUTRU3aXa8W0If2uYHNZBX
qVcRy1/h9POlAxSymKjsxRrmil1ZPsT7mUH5tlJf30MVIBqe5+UYlnwTRmyKozqpDXywxRkwE4Tr
XYQCo8kM2fTKMYmm1xBAcUrwDu2WikrTyDHB9DjS0NBjdFU+zBt6F0LFuwxOmCiSiJFoEfFlAVCQ
8ROa3Uk86aik9EkK8dNDtAMfTJub4RupA07rsGoGgSCCe/81OF38JQ4uLzSFgeTX6hr8XNPlcQa5
9mdVDs3coR0R+XvL4ZtrctzUXvLdeS4NZzA/h6fokZga+rd+IPnZDxVZRB0B91SJCMKVhe7FjW3G
Mc2wEKn4qnVSfyANKhSiid4bat/znBLTtlVJgLLaCehCV4lN52gMjxqmEc3pJf1WFzYPEEj4ydXa
Hk7s02gNhoZK7toxrxLbCABpn2H0Ppl0GPTcpMwbcYs+pCljQlixbhF3mqVeASzlvAbp3h4+hOVV
TU6Kq0UE4dkIvexV0ZlB9u+DYWAS2YY/ZCWuYqsLBlTqcJP3YReNes6n+BvlwPvLG8ET5nPXZq0/
JcbUu5w34v8t7s5Tl4fmJ3FC90NQnYju0nrRvT8O0jK/RAOo1jQoOQx93Fd+AyhPXjSUgecbiyxQ
2wsbN/vT/sRS1Lcq7Mc1k7h2A7bNC2F6rxuci5mlXCgH04Mk6Ne7FncwQAmJ6t/HmpjHcRthHC2y
07BM+7c/hWmu7kgANpOxqDl3GE5ZIS4nsewfLDqfPHP4Zcyui9lBNIbZexYbJReWkG6Cup6bhY2C
/Ri8rK4imfAUJ86DhQp6U83jiMPr9NtBhqzvPMHUax1EVGTswdlbRHrtS6qovelBMK8iPguAVYrO
r3+zngvR2GxPgg65O8gHgIk44yekL3VXv/u4OXOHWHCAYoejdVWYeshDHa80LGAXcqeZ+JshL1gV
5NaphRS/Qc+FsNwjoL8OGXXnJ9Olci2mQXFW5zxV/lJ+sRHmUSGuFvQ+xBpSMJfbcGAXvnIo8p6I
CbykiyiBcSFxB++xK+tLctCifPa3Ci66Hq17W0Uo7uGNZrDVd2viKJ9c31/Ll+rz8u92GjD9geIb
t/PfNbYDobf46gSY7jCOQKQuhFi/pM7+NS5M7HLuS54BgzToLDTMWen2JHEJw2kAHtiEtEXeXwnW
bpup5ntsJ/B3uZIb0GAa3X4jwsqiNiBwY6jDUZKRrfZ3EAyy+xqJ7SxLCZBqeJN5tI6fuSvtgE8D
dH7/bzpzhBpTMBVyj/loa13YC7OB2E515nOkP5hIF2ciSoEdZ1FxRIQZmnUm+FIDEUd3562loAZZ
baDCmHjYjKeJ55aFaKYdYvbheA7Vi01x22spif7zi3PCFrvxvP0VzAFR1GZBKkar1frZ/4h+eEnb
gjTazXqhJEB7V2e5IA78Jawd3JEa/n1FlplApGSZG1cFJLbbnabbnSYJ59CRKtYrpChZTbQ9cX9D
3cM4DEejxmI9Pq1Yiw56yf9skUjTyh1ofoI2WrB3SionrDwLQgWcPE7lZiEL+hB5FZuaAG2nbCmZ
JS1adorXsm1ZNo6IblJ7Zhevd6Vb7ivwFk63B1C10x49UZcDfdc7D4nTECEQ8ar0s+I9LJMPAEuN
beyBHoUdxJl+UXbthg/hnmM1tCAz1LJBQGPUN2KmPib6S23uszOvBSmUGQ4wyoIOUIrKm0h3S7jk
gGnDPd4FGcYH3AAUecL6jamxJac7jeedNjg6NR96VebIQsOaY+zRlXrPDgz8ilKKSmtsvXOIvYl+
3aDdBd++LdPZ9n2SlmDy3mboKwF5wH1H9ZBCPq1xOw0c34nNoog5Qoe2jqVp182hLdzBUwCWo7OH
iEOX5y6IKxhD/cSDgsWWdcyBjXDfe9xmvcocUcLA+8mMKxhCH5YK5unILwSGu3TvIDbb+R5uPly4
sRqSFWFTR6FWY+3kS3jvXqwIhYgeoV0t6ix7/Sbp7WYOctN6w08S1vg52iUdF8sLpTt3Q0kQzIWE
vQ2Zsk2bSdNKblr72B9Z8dCBrLKMNJplskLpTxnvLt0BmwQfCtK9ztnNiODCprO8v4WfTayLpOd9
XDZ2PRuk74mFG4nW/UN9+J2VTQhqTbNyIUUivZYRX1yrZydS6ZrmDOjKJnZzhM/O1mH+SGQ+3P3/
dnd2qMY3+PB1PvsxrFat6ZJ0H6rpTsnws1hcTNuXxpb5E8axs1vM59YX5sSXIWkvGdYGjHo/ravy
hbION9DXmWG/RhQhBeszv3yx2BpDo3Hxcr8+XDvcpFu8UsaM3dc8R2OfgzYVELs8178koU2+HbiQ
dV5eWXAJKCmMhLq5W5fPA436NUPgqid2R0/NtpsJny+CX05/8/IEl2d7oLdMRz5P+nByobCU9w/q
4n1f9xF7Feq17us08dtRISHG2M2klsbC7D7dB+rnbg22iWyjb6OuiQT1C9r99MEom5umxI3NfBbg
Tl4yUYoYBYsfmFmpgt8AnLlDu5tJr1IJW96dsjPEwNrlJOp7982G6+zNxDTs0/I7hec/DY6lXnAK
zfVIU2u0QI1D3aqBuMTmSlSpCWhb3sNtK2z7uC248multRlVPvJZojcfKlWfpcBerSodtngRASSl
lL52OMSZ4S4jFUtDeHFX7PRSgj1xudefD6ujOVxDmOUV1t1nwTWe8f0u2vR7VuLz6NYdKNvo02Xo
Z+/6UyLycGNfNPbT7QtVk2uY7oJLHj+eYNvnfNpEwyr2TipjduNGnS8PsqkGy3OdPmq8NuEhtYuo
/kNgjryGnRsO87Coej+DuAoqomwsEwZnhnjO77bfDCy4Lt9f2FlnGcSe5XqOTh9bOgeRWF1Wkrlq
yi8BgXuUY7pM8EjbHLG9u4k0/mGewLW86u6W84UEbB7ULw1tA6Hw5/KoWDyM8E9+TpAPZpVtyttu
cj39iFw6pN01fct7Ey6UwK/1h4QjypKsEKKDDPdGD9pPgYhA4rBSgaPRaAlu3ZgTJeE7MRSgNTav
KrfXSt0wLM4a1fLY1RlQKpR9yXpsZfOU0gg0PdjTlbllppQooeISylAecpbzXNLnhRmJ0luWQ5f3
pDJvCyQ2u+vCx4UurgSUOTaFEOQHR5PwVSxUcIn1b/c52BDP/p+6VUpopJjz4QWwVPXJ9WRYNpnf
SL5yLr+ZzsPJO3JswYMTlXOaCYGkVq0tw5aIMSAO+17L5A5P86HDYycCVVM1txR2zXOVEX0bSh8i
v6XH/mKPN/3kk22/GGPgv71kwJXn67JS7N2KiBWRTV9Pi6TEkv0dT74t+/e5zBxJnM6Ced12+CiW
Z2KxK1f+leAIf7cHrJq/h/SWF0Rv3Xj0RfbmvxR2qkclYd5Mie1ufrAp0uODxFYJX74OrDrBX2aB
rbHDGUdP4NqmK9sjKhuE5iyqsDDVDuVJusdxkRUGbKOFmyNxUCB4XDC8QYewOnrcF7M4DrHtYaSJ
qNmo4801GFnatmOg6oq51sv0xrnnu40TsE8Acza2H04GPyZG4ZKrG0okrfSvPchxwaXtRdPHdZL4
hMEYqTKxBWYkq6U7Pfa5c85iuCLptI8N+5G3+6mQr8pZooj0jxH5KLEfToMypPDLorMngSFqRRZC
giPIeSb/bPowpn0ZYR1QCL7UxDlEE4JD+L1ncd12XmYQW7VVn5c970VzEjyXkf89OBv71rgLLNIt
2yCqgyFp58w/Qh2/UyGgXkbPPwNr7SGF8/CuCbTog9Qn3Q41Kfs8Nh0H/xQU+CnJtrOJI4IA4+yh
RXTXsuSxRTl/1EkOZkL4oTIdYuevDZgDpuLvHEdy2DAhvS8hz+4VtcYU4AyLZzkT7qgUKyiHZN86
kcShg95IPOdlBLeTGv9Yp9wIOmMoJYCebPG52p5gby3LWxUK3D2dAsqzRCf9u2YlAe+2emNFnaEC
thSRquiNVO1zpj/L9NeXJ2LAqsnt9O9aujFBNzJKi+ZsAFtikpAXCi6fFvFxjlLnHMlleW6Ai8RV
EF59/wLOZrbrMZb3Zf6ZyaB8kG27rxB9+1wT9m/gIefVteWmisCq2iCCiFmIrOzFV4+kN12IEjeq
Jekce2qlDUauJO4FPZZZgroyWggP0nsfQHi14F6kG4cynGQX72GWERF1sL/c7OwY5Sk0Qo6CAxBM
DU5pnD4M/TGJjsXoeVsP1badCtoDY8wOP96nvjKCF4kn42qq5CeP/d30RwczuzKkoone+NK0petg
LpjaIpxheDXvvtv/v84w07A7WPtcb4tfW0MHCR5qJorJTs3vRPNz9d/omfcGlWgbbPhqZCZvewh4
9Z7E0dMyKQUPe7S5G1Y8gw8Sj09hAc7uOcZFCbVDIt8Nv+aa3SYON5JnErJbTZ4JYKeMLcKjH/LR
kAw6KUGiWoMPY7gHRzKITLyofiofxdxzq0ZE0cZR9OAFQcOw7x7SsyB4psYZABuGQJKuqXHWX9+r
UeEKPDThXavQy2SaXA2w7nSu2XhI9BDayQ1MeM8BIAGCaHX5tgqvQXVK8loxdB+Mp9/Lfoyj+9ui
73SwAhV3n2LfPDi4Fu0UHLTCvSMFGJDJ5RPwvbWa6dvlgyLG/3KMt+CzfhQVeT8KxuYAqS1v+jqF
rscu/CVvvxTBBUEODdgwUGflLBmV4eiCvxD+qbParWHa/NoO5uQlrPkExRNH1AXriu6TnDqwtaCK
x9IXVbmBG+wbuiyHiDwIC6utisJuzENoIO729O5xYES4RUYcthbIQQUGHRIY/JAWWY9T08ivnylP
GGC9Lhegvskd/CuvCz2afhxjoupLesLW1DfXC4sJk3YTdVojx/TScIQgdKWRTwhm5bhSillkLlIT
33/pG59rvVBV5rC4jpUSnubmw1jWLiX3VprqT3m9mnym1ITN5rr8lxjQ5LJRHFyDw9lt/JX4kEsq
pQa67ovxRH3V2HKQ8rG4AJIWQqHOT+Cs9qIrUWa0RkLHtmgcZfxIiAvK0MImiYkm4OTvyBytUjCO
ZDkIqZp30u058kOmP6HkPOQi2HXn7fawXDjgzsFBk6QoPEwZiR70Yn8iWVmsotKM3gEGWx0ST2lI
mvaT+SBkVplZdSL/Y0A9OFrkYnxjbE61z+rxpKx7Z6pmXl6caDenXlAplwenzAmRKlrgKHPkWTmf
uwbRR29t9PxBXKIWj4e0D3RJjUgW02KTzJHm3n3y14aRtncpk7jQxFhGXF7ogN++7UzvmA5d5pbj
60r2J3THWsqHap6bXlqCAo9pFIcQ+s6u7h8M0r4BDhNyrUHkWY7tNYO5GKHgFF6H3VQ7gYpel0ct
09D95p2PvRkONxXLQNyUivIYfLqrLguBVWFt2xk7A73yL7jHZiyQzY4AQP2XwsoYeFrGse2/e0tp
n5fFOzQ+NnJCEBNz4q53x8jjJpnrDVTI1p87j9JNhoQ64lQYZRIrkjJ0iQIMPTRBu5v6o65Qd3yb
KH7j2u3+QO6N7aarh0+a6Dph1FgH1S3XZts6HC9c+aeJK3HuN5ppwahbUNmmnkA3wRMxc27+hiNN
CZ7dmZCO8o7KjO4Ov7P7sTnLwPS7EDjC/iMVisCwt96R4nE9ZNNr5ZsrtBS9hULt9bC50ORrIATo
SE9kHhX1MOOo3QdW7lXHsoLZSVqyBz9j7nr7oB03OauAgov6Z9BjAEuS8Ab+VvQyxqhrabUNxasq
WASB5B3noyPEOtQOQK3ZryVn5N+GZbOJ29RS1OAu7hkmVY0Er9g8Oz8d1OAAuD3i3jTlSQyoVrr9
ZbszvxoxwOI3ZV5lSSAzuNTk1AHB1FXOWA974wv9UMdeqO3feKR9X7mJ7qN8PgNZMxPdk1ii65i8
/OGOtYsCiJJd2HGsIl2fNj+9NaBXfm3eO0lBf44tBIWwHQQrbcLMjtUCZsjSOvaoA2dTJFvSDV/F
XcRs7aeuqoePV4AFMdDtG0Y6EwV4dtUe0yyAaauM60c7WIH1NGVCtwlv2+HWQ19sFoUdRAqSoF9g
kf7BOTKY780dFIFDvA+MVSoaqRgvvzy2Rw53djX2JgE83+UvkHiawvDVqk3+vV1FKgV9vlWo2iuE
1ESSjoacrVSA+CO+6wqzbRCy7ffqLxov1B8kXwnF5fikmkCg/TG7YcH7x9lytnsviirU2dpswYHf
JytkMSLIoYT4GO7gSQrSgPMP3P1WzPfIRLJDctr3eamATRtyLTOnAay953UqMqVotUPbHIUlz2jx
hSnpdlhKDLlg5iZLFdJ7hM+8f8xNP9DcWi9OICmh3V3HKHXgnbyBgLvaIRQnfwmTu7RW16s82bzb
00azvOAF1Bz8Xx8n9DSPRzH0wEdsk03yqSd/kMWBa6d1IWGpPL3nGDMavbe1aWr/x/g5SH4YmP+M
yT3FrhDwOrXieRAXUHKWX7wXx3quI1/HROW3QYgd45JqCo12VYBJMmqk35HwLTBXx/ZoM+aolmjc
Uj5DaQWCAzAnfu4bj5OUWnlGFpOvy9gg7CC3cwjKAr7k6lNY87b6aawdBYbkoqVgStHy8uk8P9rv
AnHC4NbvD1A2T02gPCApmNpUlYb2VNWoYws0Q8ApFfPx08r0CDslQ64L8Et5M0TAPyAsDIiNoruc
k+HuFZv5FG8qyB0/8mWj541WTnLhuBAo7oxP3V8jamGaiebVtVX37XpjGTClpHyDKg0m0gZXp1IT
02cLLl9VchYMGGnTCYmlbupc5XFiIaRfig7Lnd7BdQEnY2SrbnrNrKoV9K9nDB3NmzIO5Iy7EAkn
HFQuDmgUJZUdcaR7Vcm+cwcboSwDC7mguLIYZ6TKRU2XyHAEtXOLiTMi7aqN2H4gLweoyImoIHQd
8cdVyQqRI2A3UJIZP/SzKOA+9Kz7wkFy4TZjejJcqj2hAHpGl7tpkwBVA9gnwdlrii5qWqUjYMHp
Js0f/zy+BrE8wyyOnixrxP5hnIoK2fR8cQgPV29dAhK5cJYaJ7knh3ZJrfUDB34PJ8s0Yfhxf0BL
Bl1CyIW4og2sDZnrkAczi/0fpgK/karZkkLTToR7MMU7/PVkKVPSJXlutj7ggaOTKN6g0upKoJL0
5z6Nn1qQTqMPV9zQC9zbMCP/vamHzk0dPSnMajLAeips8Ji/tnwS2dMWOqZPDy5kCAu7TAkpFcP5
SORg6/WqzEVyrk0nG44NB2JHGZpJbPTuj2+9KK/QeNcv2GzOWXWktExZ1bwkikeSfKs5GWMWGTwh
fN6irmHXGeq+/SqiWsJATAh5CI5QMALdH23uT4Ox6NtkX5KM0zbEivqUNZb1gi2/bh5BUDKyaKTu
b3Kk1OLqrV4OxWS/3AteQkAvfSkMxH8cFIz07zg1FXowZZm1nMCuvvmLXQ9ncihrAOtENNNEWJk5
1oRot1hGDhDxnP4dq/VVasRereXOqdboIhZ9J+adJPjHdHQtv4Hw30W7DMaCXsfhWLMZFRQXfp6b
bOBDJJN2flh5gudq9oGp2XDHv+t4cM2MH9fZibqKjZH75RUwMtbkzT9laF9u0dZRnPbw2YAoYedI
n8x/zG+mLdQ6KHQBtfCU0yCkmnJOfGi2sQfH9Zfc2EeRl5jvmJS13UqMAYeztRjRUH04yLa9Oecn
FSELUUKZbhHeGJeI9Qbx+8wPeWpX1kPC18y+JSfgsp1vy7iwdc5oUuiEiPIp2VbUNOd6/IW+5ezk
Zz4uRfqVKEH6FGnOF25XmA698NPfKiZpzZVLbOsw2jEBQ4eUlzEWo9bGoJkUW73+yM/75tS4IR2S
+9C2xdtlok2As3raOg+QamvgL/ZdBojOIlI4FzuVTr5knJpHil/prTcAGVr/GnBooQxYIzOONqKv
IKUWrsBSya/X3+3CNmSP4hGNMxkpnp8ATfDaI6LqlQAZ63Hc1lRicBGk2yp9oDB1mh4ZQWxrPPo9
1TZfERs157I14UeqonbB9ZnLnhWgrt4BStESKQ9l/Te8N29rafP6PpB2twWaflZ7qDNnjaDHBhE7
Jx2/OTsvK8/OlIJpBvoVQKbnEOSx+NWF9sBlzjaXw2opd+/PhHnMN4RLGnwxdNRWIVghfW1TBZ9M
rEuGsAMZb1S8aua64EDzh5gLXeIA9lk5j9M0kSq2zqPy9M9ZQ0FnFBQFxe3d1P/EUIRvX30y8N1B
71obKg8ZZmO5xopSnMCwujpooGoDHf1XiMrNaJl/OOeev65DPGHL/k0CwPPgqepKe+A7Us0JNPw+
T1NSj4646c4q99reipQL38+/VPlVCY5iB+jaTrRBuL+Ye17LmL0IrzroJq1wIcNfyJtKyaeYkx5Q
3Jaoh0na3besv398vThg/Y8xzgrwyGceFgS5wuWRHBi54iXdhJ2ko8v31Oa/6DdytRrJKHen7h4P
gQNrN+Qa/RLA6fAQTpFAhIlEkKZoP4oNo3z+yj0Ee8nfwwWflBAmip1jXwy5icyPRV/wPyBwMYqx
2rfO30UlULzu4v+jN6d/lv2pDS9csl5uJRfjtHN8XYppMcIDDkAacGyv6rpMqhSiBnFtUgfTbUQg
mYvETMRtmp+jW/HFAiGcGXZtoHZ2COnn0KoVqBcnVDKjIlycZMZ3rBq38nIlCixf2fPMQXvDAk3c
ExkEaUDkg1R6b7TAktGEoRNLtr40r3dMVGSFhGU2OGpHx03U3lZudzyZYw3oH3tC+J5ztdubxyne
vg5/bOi2Uhf+jJQZi2kjrw9rQzubaE5l/QbrzndrHjnxWWYVAKlTPX9jKcaouJM+DMw13/4EhvlH
FiQWPX0q4vAzM1IgGtcW5lQuoNGKQC6WDCsQWUoClTpxEUdGBgvMoIAzcWIYJnXkbytbCXPzkyTv
1/ogtCDFwNwD+Mgbi6BQZ8Mkuhmczq5cvim3IheRO2Ly9A5c4a8hpMTgO4YCwyKKnBI+fdg+NQPt
YtSv9LyDYhIqSiDo697VNFEXE4kCrStibRZOP7O8/qzkakZSrcIXyKlhiSvOF0d/kNw4lrvCpW5O
g4p3+hgdiRuFOgWx0x6FwKzh7kzT0j2mGt1fEeJK2yTMSt5I3uDpmlmgo0onETrQqQ05oqGAFBPV
JDN4o4RjbzzRRBdKxi8vRl6FtxpKq3eVqG2ac7sJOXMfVJ5hTKBmjYeSOwLvi2Lq0z/TfHLMXytT
BEeE1AGy5NQ3UmICSlVWIcmiyqT0fTUSUheEC3nR4qKOb8WLvmtKbV/8t5ysTZmS16Ff2glFWktk
Kq2OGRvYsJydVKAopohEAaz2DQ+JcRnG3kcfp+zP2gE95KQ4iKlgMqPH3AZbDjVkHDgO9CVx4O0j
K5QmO4wVOzREGBL8vJ8WNaa9+Qs/0uqhzffHOUJXFgurcwRFpVVYv7XwInkj4L09oDm212Up1JaZ
8iWPIk1b8olI/1TOkEXhznvSX7xNSqGixdoaKg55QSN6SIeVvoVgz5yhkfTVF2Hbj2GQA46N5Xbb
mW/BnLcOuXI9pPooS0+vtxCbfdBLJ1Bjl1rzW9tCzwn97ZzEq/wqZRwprra1xYIzMN7Wr+eA+NXq
BxqZj1DOf0FlZoSweSDXQeQT8dn+OsdB7w9V1B0at/VP8OTdCHX/kEQSvIWfvt3k+rAv/QbXF2xu
Ll5lCNpiLxJbKitSBGl4xtuBWnlRuvNSC78HO4t+WMRw7PbOLQtm8ThmOyGwZhzKfu/96X2FXVua
nCXHROcx1zREUez1lh1guJzW0let5ZSQFhHKT288VNOKk1W1T7pH0vGuDPogWQnH2mNN+i3+jsyp
ZnInnalreSQtuwTghOShobciulzrPCzcTvJZe7qJkGSjcH69q6X80c50cVyIX3tZY+RsCFBxs24b
eyXg1XoLsoy58VKfQOe75puMqHu58khMIKH/z52tjYNEU+8z2Eyl4Lk81v8bGyhj3PMcHnt3QHK7
AZff9F1MCMKhHqBuipclszn5hv6t87cJHzVSZ0gUxp2U/NKSjDDdFrceVLnM6gpii0yT3uapYlZ1
3WemNS8sb2K9wZS2e1QihQ3XmLlAxHrw3ZfYPWZurmb4czpakmoXIZcHqkdc6mNh8e2ewI/CEkkc
UjETpjvtmU4avXcw1g89BcnhMRc510o5ZJYHtO2wJdmyPSsiD7TNTWkBr3QhoVMa07Rq25IFij/i
7ACaiaHEwP3f5PwbqibQbdZl3PaqdRVMDpFTnT9l9tgfwV9WqR552vgekzKqHQ62I1/+1tCWS0Ct
AHSutMNldOMS9oB6FRu61i/+8Vs6omv/PDOMedfhpuU8rObq+r1MLRYYQslAZhVHjuV5ba6N+gQ0
mT+vuPjSNvBeVuh/TpogV2GxZaCCiJjz/A24aySIp5Ulen1nH1SKPg9ZkKdsIbTar9YUA9KGzGBQ
DgNDHe+vVWWXMIXYzpxqvrpAmKGAROrrbWChfRG7aXZnRrL1fzjsMf8SoGPtQhrw1jflh/wRmmX3
pU3qBtfRauDl1yaCPrTV7zTXYS2abucfDKTPaWRrse8FgOzukRIJn9mAGiIyx7Y+wX1nWVg5TKYH
TvkLaDyUPZMw6HIkqU/VCKnJnWchQRmq1I/8+4L2HYMt4jfTyjMlqMoLtXy3Ecb6wgHcdAp8yeLD
Df59Ro/85hZ5JfCiCeMKJyi02Fr4hZWWZi5PFe0QMpAKVd9XEkYiY1C60QHkJ8ftroSmlN7XDOaO
ebWEx11mrUI8YTrtF5abgqi7tPqRobGZ/+p7ufETt7x9WTuE3fOqhCTWlq+G/eUZ6lzgGubfEfM6
z/6UZgo0hO4hy5y6K4X4+b7m8sQJITOl9sgOesTDG3scWF6aZKwBY5ralYQMv5SOJw6VlhF9uUZD
dcZQR66HxpVKrkb+aUcDu914bGnGg+axiL/9HDT0QlQLRiSq4yjwaHR8aRiQ/sgR9z4Xy5k9AAvy
UhYjotie56xYj3NXY9bDQMKUsiu8qJ/+RoovGLxgwY7YJy7rIf9xMSbOY8WkJUqkEAmSC2503Zxy
w2TlB54Iu++ScpSCszSSlMGqCY3C1S5MjNFsKhFhuUs1+LmbkXclZfUyk3oiQuuSOUmyqz8QrJSc
2Ynvn7NGsE4IE6hZOS3oyYB06rO++sny81IcgynPIpLYEqJ+ur6FwDqRXaFSZbWO6/B1vw33WE57
2JcCAlp7x/pX+kDbE18m0sehZRu68Gssd1inipeQR2KbtEJcZKr7jrCVy/BRL2G2b1774WJiyTXi
zkqzyPCzqtWNgxFy67axSl48s5Le+L1K/RYoscRQWAPrddwTTMmGqtxFL1cy4efMX4nMTUM9mLdF
CR6JKpXszQEkzHDeVx0aAHdY6d5fDjiztiJJ7mp5xdgrWJbA7vXZh44LrtEUkzgNZLIIGxQSE+WE
49f13q0bGQEIBZ2UfB2eNQlKV4UW4bEgUtHfh54Gmj6fWtKCkYq0sH97sMq3JV6FtniS99rut6DG
XjQGMvzAlk788G293iiCnK0V8xgOF/LU8dUTe+3e87RdnZNHw4AtgsQj92a7KHY/2rtqPkuZhBiY
eaXTWcmDxJFr54++FTSShdDpbOLPyIo3o1M9BgkOxFyZssvLdsLN1mnzYMBDhRJmUPnY5GnJzGwd
jQuLN49242voeWFzi8TJNvUqsMUOBd18GPpF3sVPO9IKHa0Ti886cqSIdQWatbBKh5II0n1chPlI
KwW1KQ0jAOKHihd8t9+RITdFzHHCA1Ktnk7UlDOr3B61RGAv9od8kbtmpok2L96FlJ/Qc3hNebtz
bYV4CHMaJgkuvP9yWI1+A4MDcz3ctPHgqkcNX3WjXzBHoIHDyu/szKOF6UYG+gat6VuVNiNgmcwQ
9Q1jjnsdVY5PO2VewngqJWIUN7Z5OVcNoRyCTU6Yrrum//RT0ZmHBbv/pi7iPYjNBK8oqXj12Mf6
BEq4mzFKYRvRUDeStXtVjzuWYN6e0p4kLLKMTTM+4s4kzVKwrkbvI1jqVOQ9z5m8Ly1DU5dJOqVr
ZZzqLXO0xOwFbH1rztGSL5SIR2o01DLSQlR/2QEnE9whl7eN+maR8Vn+m38iUkb6MInrEdcQbnYc
lohdfFfyWrJNKS57QT703kETGjIzo19l4CLxrthFuXsBNFCpde69ouONv/7XdQsObnQRy9qj8fMA
22JQ1Rdwb3TCT+FWdn2K/Qh1a5cwHJ6UkVRayWNsx3fHuoF6evcQcmRo+ikjipdyGc5LRCFcDsv1
dQXPr+9OyIywueMCuRCLSC1s5Mx0t3Qes53Jof4a6nrBn6JifB+a3uo14KE+QzshP7MYiBGUWqc/
lXKixq07U5p3H5Np50qeYDp5XqDZbZhV0TOjnHtrnIVWjX8BjrHvepn39aaOh/4DHH4lTi2KA17G
iDlFTRCiqyEOGh73Yz21ED3liMbWOlBMWZlgYPQM0LsX37OgUvSSJV0Gwc6zZD4q7wZ7kApeNd8a
a5kdX1Vo28t3ejzKTvJUgnPq3QJs6K8aVddxFpe/pgunsJqHBABQVlEtXsIq40GOl9T1eTwLvgtR
NrdBMEaiU4WE5Jv9wrs6OFinv2zVX804mM0rQzBlrcQOQB2SKw1excvtRyhBOYW9WYSZoMbCcEHW
y/p48J1D8mh3bb1OQ/s/DqfAki7Q/d/UbZpKiKEOEvUTn/SHuabyu4T+Db3OPPMVtFNn7puVD+Qf
fUJe8+lciUTnovy7XTLlI6J+ts6gx1q+f07MTA5wDgJFNT+p9tSzSr68JDM5TdQy8GWJW5NR1Nia
MU0wTjYT56zbeAiMGegxItzk6Df75OMYg+iX5PhRyPTSRcOtu4Rqkj9upwZF+lHTtYtZAfO3oP14
kB66XL7qvOTSpkBd84wGS2wZLnUNdM6E9uDlmJnvE0FpsR0YFNYehovRsZrFC12kBK08UN2qf5J/
9leShF+X0O/jtxvaoYK/QcYpAp9BbzxSGKXtYTSh6DHUpOGrMEO4SfmjLPk4Uz68xLAFHwXOavRw
82XrxMf7hFXmP5JMNMrap+VVcpwxfU3hVUU4CHiDr5jTiImcSO+1+Vg4+yadPEKw1MLqbkGJkHmF
7HEjRU0L/QZWym8EkN9FLc6M1wtiu7OK+BEJXmZlFWLHT63cB2jQR/GaWGuFTGgrppmyb2uJZ2wr
4tbG281vN975CDatroFGGPHh+l4jg5oR4QjzQeND/Zl9xki8combx3Z8gUhROH0T+NCY57wTpXBT
vmyqMGRatC3nYwtQQ9Z4A8pWhnwDrhMuBgPOY709/MgAo5j0xyMDpaft+HAKdUk5G8VsxMUWctu3
kIQsczvR754PmMI6g6K4hD1zPr8juKH21sXd4O9BrhhND+XrnTBxyOF8+c6y/MkVY83yHNQgS44Q
xX0d8CU5+qGClWYfYNWED1LJ5vFzJhbhRLtw/qSbj7Oxygs7qT+vNft0AYO0ToleQN90HvjCiPh7
Z+OVuF8wZyEdQ1J6WmcgkMbLmcf+uJ1fYm1AEbQLjLoXYpilkeQZZ0q1PiVtDnHyhDdLaktbLGVt
YObChbC1/TFYaAjMTYEqO9NvDp4AS5jVT/mCmhCz+VhC6yKi2r7XVagzE1ablobpuk4gH8qGVpgm
JyZ2RgN0AK/9uYA5UmEx8GvivtCX/nvLoJQhCiiXZBgg3tjoyqRpJ0x68wIWxWlYWe0JxZ30nrMH
xc+mayEypvZQa6ffjnaV4PmHtbI0B7l0zEwibar6kGkyDL/i1Oy9m5m+0MAHTUFp2yi+twMmpJXb
i04lCf05U4gmp9VpfAk/7fs+IJSRXgy8uOlWbxSwAyoMZfCuKrMrvD4OPL/YOmJGvxh9X1xIGpcx
ivSKmpXCoS4uODsrUDrWk7txa66cWoZIT2sM/Y+bFXQk6msg9AwIsVOEnbh1Yi3vBE+/6KphyIG9
bsMMmi9XBkMdrG2upcRGrNSarw2sDkaBdG+9QloW56MfcR7+opD2ZyB7OlFpOFwlYfYyHo9aVK/9
ptIdW3io5h4ruC0FIQ2viVrBe6R9MWUKUQoTLM0WXROWOL1+00z6/gG+yA9V6efc+t5JD/vagZxA
yqgPKDA+wyZyFLafezZ/XZnIC/AVkyqOpeKJ2JVItoWQJw26GBdS79cbV2foTHYFQLBBhTLPhzaQ
AjaDg+1GUW1bzpdYVVA1rlAD+LNilPJo4NqBu+Zk5Xn3ND0LL+Q6yhO0ZJ8ZkrW4WthgInaxgNu1
CBxaHosXm0sUFElMupg93zqUJ8Wmn1WkvQnYMwLJ9T6neQ4KjanV9FxlPyfBkbgkeU0k4CBFdxVp
Mfzu7UqGBy2mBVBkLkFTuZchInjNqHJZpurF6jnhxDGGU0HKFx6EnrWGJ1zDftzZVJcRp3Y8vY3F
Mqv5ywZivNiwr5F/+TmvaaU4qLOgGDLGnCIrocI50EDe+3R1S7wW9iO/FWmxUWuWtAhcixostsjp
udwIlVwCOaenTwYlGrO7JSlO2IlcwzdKVFIwvqaFuyfgGJCsufTkhKqQSMBDHZOfMSZEm0q4VNbi
dWiofDyMITIiPEItp8DfcM15OsZ+dyVDYJ0NTdIbHmadhcxZNQLZRX9Wchd/+lI2nI+Jbj673K8Y
wHCosJUaBhgRacygP/N6MGCbk733Cb3nZK/swTxbDBigzdEiWF1dj/HFuhxqDv3Zk5WUgkXMRRU6
HFmUynsJhqpUOZJ1BBUXA+x/RZOuQKEEMGNBMg1Myv4M4lYb8r2eW8mQMgHbiFVOBSHNAO0PaGiN
e59aUutHnBW17QeHQB/M1NiNcae1BF13FegO0z971L8gklNsivJdQg2CoSLkveHGopaWMTHYPNBn
neAnlosNfEDMGyQXcyNaaPPlRbeg6zNgY9i3rP6KcTYj9HTf1m0m5hS3s3ZFs9028s9Dt5p24s7e
Pa4o99399OBnCvTBh1i3N8ZlhbQq0kxn5P0cdusi6xkd0AiBm++Po5pncNCUne0dRlpxueiKN+PT
Nnl2QgPzrG1To/ilQPFXvcqo4PwR63t0brLVfsFk6IvbdYNM3YWeMVHC6jqZLog4p1amnOzKWP1D
BIFm7RHfrJySTLAhwqh5cD2WCga0acYM4iqG/Qh9vlFHxNnGD4WkOzZ3GZggo5sslBI2BKI7YXSu
peJaUtjALprf11fxPXMYlmof+xUy5tmMYEpF2/AJ01TmT1gtPjCDj6rz27ulHWA0XAC88A11Fkhl
RCJqoWIo1AGOnq/r7V1/y2kioYqR+xh5jVNn6m+KBaX6w6OGks7Lv1d14VSaE8nenbseG9OtyL0O
0HWAxA8NzjQPmTvpGRuu2OKUi3IU8LgRvOuP5ppxaUocmZa6pV1laOybxT0U7MJYZFgbdXlY3APo
eai2CgfR0fA1LyP+IVXrVddzcLsstd+tb8Gz+PRw2z/h5+1sWNnj5jbFh+HL+Byl4/zdiqrH9M/p
qv/JYpiTN/YhmJsRWgTsK5V63vWCnHAwCF56jDEZa4RzzhiFy9KQRKW1SIRnafOA7a8YwKwx8CVy
G7eSsMxqk44oei08dwXFRoIcL9k7QtKd8hIZryUj8keqwOWawJlIAQBWAx7GmWxpwgTFkGCXeGlF
MWklYYk4QCD052KqQNiNx6pZGKNoYc/ajRzeguhmy5/Ws9GyTSP0Yr0Damw8QpupmSb3k+bZOdVY
hWjW9RpJmoG40/vr4fije9CxzBtCUS1UIPvO2gIF5hgXS8SU7vDkqIHEr044c19GajNpZ+zchFUf
F7jkJrWoPh59teLMdefq4T8oPTcxFKKFpZkpec74O/wSxpbPm11E+95XuXnjjYfHqYeeS1IU5pTZ
FXFSmBRz5By39g9K95FFvP/xXnsyrz5l+KAFjx7iRso22cvogqlZRh+kPuqrMcPffciBqcK43c3V
Sc/0aB0mGX9xC2M5ZkrN8CtJ6YsIWI5DkOJkGrLhNVQ+dRlU6kfWXmzn09PI6l+jHVj/czhQ28ZF
/5GW6AZEgic8PsMIZR2znHg8UmGRN2BjS2hMQC5Wtkmh14msO/7/d3O+kGpXDlIchgZPVDlFNkES
OXtgLrtkJ+OnNKDuU+pZYQIdQRrVDOAcmH+Am+K2k+Ik4GfBfVpoQaws4+ForGtbnR4P+zkQ1w0a
gLXdPfDV1F8SylTTiw4ifGz2xThic44h06uHgIBh9Cn2e0sTw5iCycsdMlE71duj/dAa+bSf4nkw
Uz31NVpChjSP80goKF/9krge62NHGU6NF+lf4BFzsXVU5MOacF6LtWcePQwR1cWVmLzetx4+ECfr
kVAmhBNHDcj8pRXEZ7u1CwUYqN3AEWnwjaK6dFjy/9IdSGlY/Uqk6cBz6PecNQhc1vjQ9SDvX/0c
I9t1koElB0JaO1OCR8IFbpPqeGSByH07XpQDSX2mggDOorqG07JQS/hfXaTurvxSNy30NnEnhnHD
iWGA4LONHx963gpeY4SxAf3mZxdkQNpMB9d1HW+7B90DLreCaF5bSUdhcc7HmZXU96n9palgaK1v
Ml7HBZ4otev4dEg2EY5gB2LfrvW8/EaB/RG0Bxa/0+ICcuntFfFb2NQnP+jXZBkfA7g8cPRIgW4Z
kw8CUs3sKQbwAxh4Pr1DdN9hxwCbooa/wm0uBWJpMdxqnzriwA0uPXH7ud4zBwHNnAuVc5jfvxGO
9eJJwz+tBja/GPwsBje2vTWjhkhhFhDv1CibsAZ6bidWbj0Dxl+quDomfNoysbDNdmXt8BRdhmX6
0i7DuibbEp/3V/wCFSdwaZ+YlnS3N4VeAI8vDmojKttwn9AcqPxN+KPup4fXi9TIPZ6Ud2+uIvC1
XHXPL8CF4ScW6/19wSXGCvPXrZPF3TbE9Xntk/ndMhfTQjUrBNLKAhqxDRAao1njbXvWhvLmSrMJ
iEd/WpHzyRi5bOQ+z8MEeIxAFLoYDuKAR2UEzwTjwoIZPG+R1CLqFCY/6rwiPQssqQPttKKPvE4D
yqxlXm8CdLdWnXjSfuO2rI5zf3yjYmmGPAgH6IOAMoDKpnjvrOn96VRFgJ0aI+DgfYkqO06Yef1a
Z6aJS6W//qenig2nyUwMrCEnLfFdKtV3AgTCMn/DtThCBjgEcytx1jYhRqRpKX6lcdDu6CmD3YYp
08hZVreJOLClpBIC3r3FU1rrqg1Eh6ja+Snpv7L/gMFNU+5z5S3PgekJX4n7AV2ND4i/uxZ+PKrO
R9JKsaVJKiE6d+xhByzMeqH+Uu8g2URfqwq6q0/+xXxt7CvfGtld5XEdVT5pIB5AZJow/JDjeeHs
ZPxgiicaaaBPezV50w2H9hkFUps/WAYZIVJclHXP+Nl+G8qDfkfciaVMf9KCqzZHRSmL4pdkgPUx
OUhY49SB6mkTEB4Rti4cy6+Zh5SGMxpwTr83mDNn/MU0EU3dpoD0ibOLB+/oRdGtOd0l3/GotABz
7NhhzoFqNuFvldUO8+VSNECfJt6ZDCspLyHiR6ReExKAOudDHBv39CdFrGPaG1R0eUF7k24eptG5
GU1vzkwcsPpJrPhUVVGnrV3bolXbAy7R4wO6F2n7ysmfSKMg2BMcguHVN6kmMTv9/PvqoykiPjkb
OSlEeQ4PffYPGr1+J5CNd5+N32p5mc+3to5bj1l1daMCAUfq+c03W+1svXxIm32bLpp7s7X8PfTv
0eJB+i7dKKE98nDNpc45lZYn2zVXQR8BvAeGZ8jc9/f+BVv+EjWwQroUl1ztAphfoDiciuXNR9Ce
Yckyi9B+wBOTV7Z1ecGAfV0a7YK8FWGik/L3Rqz63/n5QIBQxyHyUgzZ962rIVwYsVx2TvNZe/oa
zWpWwkZZK00VDJQ7RRl5atpSX5npMIOx8N43VFwKr31AL8NG0kvzsU93SbwZTu0gvKU9+PeICz/s
ewpinn5hdgWvLdU20dllASvj+N0nrZbSe9+Hzk1ePoUt7a4nGKUuqCDJh34SRhHtpBpQ2dVONQWM
99lTPZf0QCURdUzritmzOjuTePO7TTltkEXxn3qT9X2FEuQfNvZVZyAh8kH967hU4luiA+rk/BTh
THzQ2KyajgyAoglmVBI6w6sRN0iD7u9EEeuTyDlDK35gutAmOFhzF+BV5o+5TcilkXklqn98UO1A
JJYarMD4QBVTFJ0XmqTZ9Xsz8ueucOQni5cZoTAReOPRSx5U+bV0qAgNWJuJfhytQXXTsm+Nt3gH
fXaM+qnRBgrMQtkBgyHiINwzh69A51ooKb5jfGUTod2HAYiztHvH4ZRZg7QH7QV2KLoDIT+/Ci1g
EBvPPA59j4IWTQUbtnGf8m2FkJl0fcPMeckHyyKyQv28LW5P4K3ZE1gWljnN2oRvVaK+2+e++fAC
Y2OUrwDzdhjC0/lyr9vOdrdhu/CZnsGYH3KXfd5qAWFILJlqwitz1lQLnE+YqTokZMOwGojVaD1J
mqLRaywqluZnGQ7lOzYlcpQRvHJGIIvbF1QeGb7kiQceW31ACcjvq2aJ3j8k/+YfSzcswpOW2xpW
77j4vHSyEIwy09mR5CrsS8wwHHLMJhnPSpWhmIJnTxnpIr6NzQeFIBL+VhdRaCznpWebFIVlRnWR
1uN1Kwn07tEswE3TkevhKzj5aBovGG/J98IJlpQGnUHMqjsp96TAYD1vNGzBRthX0FSu3CS1Xm/M
lAanLs0RnBTsWEarb8SuQHK8b1LihSNXu/BGpD3yS0dWFkHo3dNxgn1lx6tec0e6LVwvNAOvVngW
ox6/MPVpWnRT86LA0rwilQprYHjGzIHcuAPXG7o25NdE6mBqUvW2hi80PobhBk/SxJcBrpwe6mll
J8MBNE+L96unwfP5n8b00tsC6Dgs7t9fCiPd75CGE8esdc3NjRXYnxry97sJ4C2EBSFONKxumeLh
Xs56HWgzct1ug1RnnwRDcEq4P1rHXbKG1KTnM/bn4xa9mzQp80JARM/o4LjD528nEvRu/UI8zHvT
GS1+JqsfajRyuZxrKtxAywAMt6vTMESdetQWqNh3OrFi0tX0eEAoaoQ2vpEkAa1gIsPyif1KcYkP
n9q2dXY6nroOy5vE/ZBc/eKhbgHxczLE50gSihCDAqUQZU9ZIwqsEA34Jtaucgnqf1UJNZZU4LHs
Yh1F5UJ9Uy9L7n9s+mwesOaGgFWdN9wh3DsYVAmAxzrUaneJJ//jSpUpxNpwP3vvZDC9IDTZbKP0
G9TE/WiXwQlr2PwOKtQOn6+gOjjudpiD/VS9uTbYmVJMmFcRzNCPL2cZuOABYr2RvTec9nlpfO4g
fYVUB4r6e08eA1yLIhvPK9/qd77IFiI24RlIBjDirO+cMb+o4yQ3D6svcPB5TXktvYD5MtIyDNxV
EevS/EQeduGLsihS06ubxrxv41iVQDj6ZzHNxzSkxeh7vqFWw9Y7yvIAdR4fbV8A4ogRGjK/aMvD
ZTSBtTacq9OHuVIN4jDnMKPJECx9aZoM3/n8L9sevbZJDkVyEA5gUHhbq+6rYGp5GTuniAG9UJg7
VKr+xrrxbN9sqGUfaOIzxBzzroFMv7eoymi+BVsAg7Gnz0QrpdIc+LctHka9gkYqLuvo6TJZWj+e
cuY6k/Zlw0ldS9CHvdus2avnt/IIbirDnA3sprR5dA0aTI4kTFvamZUQMNlehPIDAiuhXZibxSku
8PNVRXoiu6rsa5hjyIVv7uafUzIfpQx5UC04s2inpnIPunJbjkv/17BtMeCzmTuUC6j1WMZ/caJp
ZWBrzpNhY+xsvE3KyNfxafKvZ2ehWjZM9R/VLRQiSYziwMxdcL5Cwu8QsPCqn+VSrdKfwETuHD5h
5IuaBGxUGt0tKRzBIbXk0s3Jgt38KaN6OKsDXUpBIgp9j9Is0q25AzUbA+J9tOeN6lAR7OiznZ2k
v2FMYWZ4Xy1/hC4+khR/KWzEGXLwKUk5gimsrS8k8QkXN7ETdLlBmv13nZYZCWs9AmJhLCRgVX34
1fqC3aIc1fFMXxlG/xKpgrTf52/5b8mi3P8czJO0VVLHGaaCL3seA+UwAhP0XCIEEJAxkRCjZrmZ
uM3fOkE6yXRxjK2icBu116fONrtPY8LkPxf2Bx/ia7s9XBmT2hGiz+eyEiwZsAD19+/Nhz4y3lqZ
V+xGtM6HIMfNCeovbvCi2efg3ADnRzRU9q/oAiniU7pvZIMPHOUWaNan762Amqp6O5bDxO3zGh4E
fcot9aAwUG1/DR6RB2C3E58xqrXZ6qdzaFU5VOJqxdD4vE2ictDoWgoOBKOBt8irgx0o2v6yVGSo
FyQRFGwidius2eegt0n0Bt4D7LaP/A5cRP81jJs1Zk/rC5iPbJ3eGdukNy8h3hcAFb54CBl/m5WT
lywWDFAE/1/KMXbO0NaJhTbyKNlqnZcBo6ZNOHLyZlXdwo+xSHSZqBkUM716En2eQLBp9OZa3s7L
sFXxs1XU39WW301j8Ncn3dZ598+SS9s0KBIcowyGj/27ZkOdpqypLvY8ewB5Uci6OTajkbYaxPN1
adsSa2Me4IfE7RZgfghv/P7wbTDxdnitKJHkPUcwwvVQWn1bXw++b2wYAI/ycrHwjdky2fh8+1fI
NyYGDItEHzrKE6Su81M4XqKvSVcNmhFURVtWcRHUcZqPuGENK2+y+RLaj0UUFlxZW0toIBRJoI3L
xEbgN8s8pY/+18331x2R8DpTt3+dYMZIPu5+K2B4VkQPkDZ+ACLJv9Qeabc1gz9vxh9iH7AlGaux
sDAwdtU0JV598JR1YOJhSSeQHYiM3Ltds5tILaRNJzu3+mrnNZrr0WCPGCODfvobuXPwU/5022oj
MgwnxJB8n/I5cLWJByu/g55P0A3ce2QF/lstHMkR/OCU7pk1P7LgGonG7lQPDrv/cKN9eEc0KHYF
dsYvNcJtwpUcJtNMSm3SvhbbRRCLXWq39/IpMhN1ROBUb2lnBYxaQJWHJtAS4YW6adSrkJ5j+RE2
TFh0BS4TXTXLWnaOywwUUjlM+h9fU5VrYB6vXTJGhhltYLnyEuxEEa1BvKNZtjZS+dhimtQiuSpq
yRX6l/4aBePq6gRMEPNK0DuClGZJXbJ67SYNA4427PAded+pFxTHKcdeW5xBBG3lEz85fMJll54B
ms+/jJIxeSmrXwJ4wIoKG8r6fcYSNr/J5b0Z9evtx2ZpNfCZBOcY2hgC3UwvB/KA0cphyT1DbN2C
g3nNcZh62v0VJ5PR2U1yqMyONZaFwQlTStRvBWxaV3QK1Pc6Jo6E9DOBQ8HgugiIxPxcttWQ9lzz
2VMGyxOMF+Bj4YtkC8aDwNfloRUbPd/r3L4Pyc/kJTI6I0B2h5Nl/A5d9xGmB/bspXbIf/jdFSwm
OO7P9bZg8h7o7xG0Wy0AUN8JG2vMGs516AASzrJMiE2A8l58MfQ0NOvlJW0AhDPnNJyeCDpoxoRZ
3cubfltAV2ut62Kd0OtWrO0NJbR+6rAadmWaCBwGzDsa/RNYBLkX1L5P7JK9KOq0gRE1PSpoExot
iyYNb7hXaRubfd4Sqa8RuJATrBN8n4RPa2br4391H74VVcDcLhkiuGPFpgpMnPuz/VFOyF4wYOXo
OcDLAfRw/uqpDqQUKutP1xh1rdtACqH2u9MtlWXmielOfhMRuGcZb9NDAwNX9HPrND6THtAgIdK6
hMU7tYsPmzaxtYT7PVqMLzGYr1oMLdSdWQy7RBMbc8vKaeIoriqe2Yw6wZKrOEbRFO5e6hdUHNNp
VlJC5coaJIT/OOZXVSiErOhUC0cTt6sQiXUNDmD/V2gVQnZWjMBCziB3SC9toaZE/JL3Qz9HXBua
fioRzoG6WVidj+ojINuoO4hSfLwGwLLZLRV0PiE4jSq/bT1dAnUdYWb+h4YaNt6QIFs3Nk740UcQ
YtJoNKEOCXPH8KnZFi9K9VL4HL46ALFxmVLnVh3EmkZgJbPPJCXBc0gB0QS9gat5azmG6NtMXE3J
iJsDCCp42KbZNsh98k/Qq+aLOFcDPxblazxgwdDCDyuFIvgZH3Rw7djCdt60lzZSF/1xuNC0TCZu
Nm0IlvW+VZOfOGlD+OSbEetfOBa5gZx4zGMp2Ji2l37k5EiTxNRMt81Jp3taT2FIN1ffm6AZOLSA
NNXg4wBmQn2DEVa3FbJx5PZ8HK9ptelD2thXMi1fheJvHB+lfXND35eXNTHPJOeMIEjdruFPV2TH
9Q47MPlQ5N+dWeSzDg8nbWaQTHesrr6EC+/C6vHC9x0HaVoGfmjQgymvZ0V1JCVpH4dAezviUoCT
/XOsSDisW2fatloAr5ITPjUqexv7c3r4a5NPivO59HnLo50eq939tmH6kAYJvtHfk2qyYg3uIdbd
nXjbW/7C2HoWmnEwwYxgW5bdzyk7184djlZN9aLCYGYXC1yUTzf+SRt+g/N3Ok9yZM22MSYD5X89
bM34JfxcATIdFuzL2JA4g/ZLcSzuDovIFcz7V1mV3dj8vRm2ePn37ehz7+Yg899nKr/LoK/SV/mE
2CzxrRkKAx8l/gZqyOTRfC6RrHLIAoIuJ4KlBNLrZsU+xKToVDpPXjmCD+4SOvy44kBRLh2hqgzI
OkLmUJf9L6UruUv15Bf4HxR4JkAZZZXjxTFRADsM7RVRF3aXkvDmqcg0+I/LfWK1a1Dy/dyWZbWG
oH7MGgDJFm2XI9fiYCr2dmJA4llQMGEXwkAH3FiP9+2uyOtU3+IhL2Ar9f5gEym7FwIaTMamRT99
MpW8MAukCmnVGs/LySbMOo+kTnwAsVqxIiXyxgvK9zQjzXrJqYRQYXodrZp+KR3HJpvLcvGReAbX
k4C6Zbl3UTiEwZrVl7PndN2w9PuSjup3Ihqaq4BS7JpGImlx8ijYWl73+9yqNaKOVcGgKxSjMGS0
G7j8x7bCwM4YY0fyZ7crTH29STM7RGMuciJ6GkVaT1vXXxph78bVtU3Eq5pVGJExufocngkbN/Yj
aA9q+fO8kK3iFzO3v3UKdDx9XMK6mo5fzIOEh6/fYc4jcuM9qs4F2R/bEjlNfZ9GdA4S0dqH83Py
Zrzij+ijascpxfij67WioVuQUNTe3mNAXIZ0azolRUOq6/+joolX6BYL/Pmdf2fEd+2kXHjsC1V9
Zo9JK3sV9VF54IEKu0/ZTD+kGWhKz/tljAcyo3eikkD6T3Uci5JA+s+bXDTFfDFsdIVxnIQAFe19
hW+eXwx3wqtjT68EXol+fIWywvCAvUt17k1KF8wBSQ43jbqjfmRjLPrFuosPIdZ29NYb1fCItKFI
pZiXT3MTlfuoyYsAQ/0OcG/OIx30qhCsgb+6civpszZAAwKainuckN9TwPFeS6mEmTXFrxZRr1h4
ONBUU4bVxLZZh+eKxENU8oQHl50x2yllcJvXbYRGjAQcWW1jSAKwprofN+UL9knmilVPF3sygsn5
TfbRtgnao3pDUfbbJw3j3Af31S1NERI+aD45/eQyXAT3OPpi0HvA2OsX2GA+9AqWAocok6S2R/Pk
DoShbQC1oDaUHXHdnsLGy/Dch0AzfHMG7bbw86A0Ce3G3q9fiiloTvpwGIb9DSu8veq6tniwN/T3
tLJYittfB5rsra7xmL36NItwm6ApokGjjdJ7WNgtI/TF2wfmPG3S/eDC0mrbtx6jT0DaHQ6q30Ic
+x0Ir/EQ0mk3nOu9itSezbh7mlKXHHjXqHbr/mQuAF/zqJvfi+3TtalooqP2a9fAWstjHFcj+4e8
hDEvtTUwVcvVEGB7AfH12toNULRz1FI5cFqZC72FfJw06//tPlMcZTEMxb9+HLAmHb1ygHky5q1v
Q3wGzlusrnLWNd2phjjVy7JHWsIjGWeTudzNz4Pz89X2uGGPzk2dpCn9AZ4v3K/yVlsTlDTdJuRD
KCBaZmB4rO0HpqKVzE6CDpYDfng2H4brK/FrQk6rEQZOe6DvIqxeCs3FgbRK5jp/PTQQSpZOsD+V
3FLLTHeHP8ETmfhJ+FUwi+uGzU6GdPAlKqJt4rHpsIGnH57v1vYQJPpzRno1OLd23O/OHCENIJ/f
jB8c9L/qPCmREQS2o9l8SFUfCQlmmUo4XbnJpFMDtW/k7h6mt13n/w21MvXeq9cBPJLpzIX4Ktg1
i8kdDThd0AKyI/rGvlLEgZ6uP6SJ2fhhHdgPvnHJd1Z5sUu3jRBozLLg2gnYLs3aH4wGtsH/nz0x
A+nBTNLRSkba6624nKyGX4BSyhmk6TYyUldm5DC71zfvS07UA7PYnlvXuRAOgpGMxhmOEiaPDwMm
eypEh6ibKodkbaQJIifH0xvWj1QrVzPuz81Q2Q6K4TXVBODfcBeL8AM2YD/teu8y5En2wi/+ScC9
CYJWV8glCerrW1/5qs3qlNPHAEc0tsUtVywbrfkC0kIBSV+mpSta6DWnd7cVW+wwvVkv81DzqWSu
rBRZ/GqUwO0v6jJ/rnRzGy6UXM82CtgW7xTl4Io6T2qL5zgTU65EqPg9VPlTlri7lkAIsA4EaDis
QxEsVA2mceLzAm2du5Go9JJKKa/9hruhABOE2XJnIrRWmdGfoB8JFgi+3mn3JO6E7netIPIOGjqy
38f8XURV/ZhAqdIb2K0DipkWWGVGHh2TWiFaFZDgdiDKhS0vULRG1nKao3atbfXjVWtDFi+jREmZ
QqF3hn/j4nzQ32ksNhZqrZ27CcU8Rn0WoxNqdoFKFVsuWBQRmETcWht2RaLATglgPDMGGb5Rvmeq
TVanmp6gBFyARmerChEaoHHF+TlJHbzO7ERcxqRf5HI8qAHM4JctpZCCKm9+DOsAjXdSqEa2ptiI
C6Dx0TdirQP8yXHYtpqpKWY1jJI2B0ldEZJhPvigo4za0ixaOHb7NNEIdG3zenQt2N1Fl3T4x4Ph
sk456vZS3rasBloF/ZLmzzcOvsSEnBGzQO/GBhxmjadEPFCwFTQn2+aN8DUDI5NAL7OBKLZzOaoP
JfOitJlUnDbSo64Be26dw1KQ+jQfYsaaQPIaZfwbE/VbM9lHFit6/gLlpK6DE8aem5BBiB9W0cJU
YvMKVx4ImRRRpZzqmTxFhEZc+EGrQcyeSmgDL6hB6KnuYc5RQv7kFfe7vm9xKRAyv23ldiScOBgJ
W6dWxiLtI40VzSiOfS69MytuRGg7vtZ/WTgF+ET4E4uS55C41LfwMhfDvsErbo4Uxn3C8Ln34yYa
KaeRaAfOenXkiqKUNFcAmS0SlK9KPimB0GxMwPSQOBnieS7anmdIMd5D7DllJK+ky73ncMQJqMbH
SY5c/39GdQRijuiFxT/Van/6LjP3VIxRpYDRELZgeYPQm8l5MT8kwlrzxOoVbwoAfCe7sAZ/3wsb
LrSjl4xRefafBRbyNRNoXpQQUm00PELx5wlcl2Quc6v1bhbR8vXlHI6FUE454VaCSGVFEpOPcM0j
HdfEKRR6l6G7cV39Z3cBCrom5/4QFgg5gQR3zQBpLLHRq7vJYZPSE2s9jkymY8fQDwNSSB+qRzfl
bMGhTAfvGJi8Ts0sWRs0ZNHYJ4JFf9ILKqX1Vdsi9gz1VqHZ+f4ZiKqiuHaDrRdwu9Ote7lxbHek
/UUme3vj2+DJ6d9cYxuGywkmDCXuYsfAlAeBbt+IgnS2DysaIaHAklArU+LeThQ+RU3SCXAgc46p
SBcfAa6OKUP2wAU5L1NwGSUM/AmeINpAfBnBRoJzRswVC2bvzxtjl5LHrfqn0Gbvdg1Z6PHaTEJ4
mluHMiMLDgQAxsMEc4qIKCodhULHjtb3M2jaQRvAXyZjN56+IOMWX/hQctuoOkur3WQnbrSxRYrJ
ds6ZGMGkn++vxeL79ecj1hUJ+U8ZJ/lqU9BuEydViEVqcqvY9fh75IDGCIyxlNwttBbXi7MpCQKE
m0FRJ7eLdcxtVx4myO1nOq4QCRodXWrLilE6IK1UrRmhMbiEOmg9e+fpEmRZNQyFYTpEsArP7MzI
Mx5u0s4eudPjALzis0RWqHCHabUX9+7qnmY9ebsFC2afFbSBDRRzl9aQey1KKvw3C9+3X0C+WWhm
BuIZi/FrsqcmLS1xBgbkQM6Ip7e7Yq8wjSxHkNrw/zbGzaSfp3sGQxWGLYZFEY/C/bbKhoPnlfl9
dQ1hDukiNPgxE5YF0AQs6vLmeu67YhUI7oc1h/pcicOQE5CsLEIfg9vJQYlyTaHNLCv12i2ZqWgm
mE0c82Ds1taKllKaSnYg4he77BKuHq+eIEEFSJyaNT5naGJ7nlrHqDhyuGuyiZjKD9jYfvbrJ1/Q
0mnmTEDNlPjF02zO2LgJm1fp/D5lox2rlLy6/oMeRdkZ7N+QDKmn/2F1V31LYHS2BXhFKTqqRuRj
8HEEZxd+HgHSlI36KDb3rq+sjHPOIkzFNcAvxAJ6+AND0kSiwUhQruJ8GR32QGdWOoxiTvK13qjs
8DQZbtTX92jKnKiUaGpJaHdN11hUGvJnyQDgWm/uyjd+RW0hHpoLP3JdiTYPRlr4oga1YaTpmGuQ
zqggTDS9CE6FoCWOGJrdoijlg3FikC/KiGGh7/aXC33D4GtqGG0dV4OOdD7xf4caScaIpTPzXakI
nxQr81esq1d0CdTWASS6F/t6mwnprdtocwFDOtGJr4rzpvTmLkNlul5TTr8umXiA9MCZF6/wdntx
6EZJnZg6kcBAjrbfoNWKQe0IMGAg7WfWHO9owHZxLp9NY4jjm224EPeWjE/TJQWrocdsafXZMmJQ
zhbGhQSLsx8HUt/9ahGkYY49sVRFuTtih98MuCoOxT4BQVSbCI8FfpRWzuj4/yNA9iOaOOBcTnaS
6dii/R3+7yfvcBvV0TCsRuHinjR4TovEqPrRR05kMNtWmgOkz9K5mshDVgk8EitRvlohzgIaH8Vn
G+MUBJjW8+wZIW7k72vm37BdjoBP+9BB6R+9WYWYpmGbG4jNOlYQx5B01ylldIX9tgCR1lGMW1JU
8xhP31koAEsh3OXdsjkC8GUvwFoU1SW0IWU2e1DDgL3btDk7BRDnU44mMSt46w1PSW8fwPWausQs
toVGxT0SSR7Hd6slmtLZtW1/wW3hax/HQReUHZ90WyQ+e4q/aIOdotpKaYVTD7wVgjObPdzR4/yp
vaBMnUjvWYA8EoRzd6izUHIzKcViP4kyxK61RvhuwDlC7yBDTabV9gTD41VsnYPNaGxyNfeLqCaF
ke8oDzTpm2242nPMHlFDHrZh/BMv9KasI08uMyV5RnWvw5407Q0tm9p3v3Ns94g903rK/REaE79r
YdJgf1PPJFEQXSHT0hyNEZ5sQ2ytWPod/Bo9x7Hkk0SDMaX78XhNRrd+7XKuBOIWmYZtk68998Ke
+kRRK0YsCB4UPkK3WcU3aM9lHKe90jRP7xWZ9XWviIbw5Lwewshkiij0g6es8lEOfSBXqQ8rdqZl
AJgQJutS2jX9jE5mVbCcXr9MFORpCqY6trg1zR8IAFokcF/yc9IO8zMahC+LmvH5Jme509Rfz+mv
+huHBw03KMeSy2IK6QyX+8DB9KXWSxnl5bMQ8rI3WeTw/MyIn4c5LWKpWsGQ4W1+ExgYSoir9MvH
WOZPQjEiow+xAkFUiEUZ0iLJOS5omImdL2aEzCDWlRcBLAPM1Whz9Vt82YgRjMKwVSDsvt4CvGW9
f86kLDko8+Npcit+yzsveD5yT2r9c4S8ZL61awOucWddgKwRq/shVDmjdZKfaWmZNXwPRlcWdqaP
RfRerFvjt1cQQNNM100VI8WWR7NnFbRQaj2mrcmnr++zty0zq2Zt6l2/WKRrxj8GfN0/mm7qwIpb
2E2P8/sFNd2UYFxGcRPIZh1HwaSzR3CT1Cp9Cmb+cwnUaGiu5tJom9N5ng4O22F6CyTKHAWbBH+S
NvBNuM64WIxs+qgumGJIX82j2CF8Pmt/uW21HjbmDrTqgUe2hMorheSBHIt9PsWSoFDHdQaJq2S0
uNDYAqaHiwb96bIXo7zRYxmg2UCP/fT/5AG5oGKZYDx50L2JQ4VGfg8IeJyjsWvZysQMbMOGCPhe
AN+T7I+bxIFtaVbnNytxy8PImfBwn/by5IodlN/zAaokdqJecGvDg/6SlaP/JMjH6nc8bqmfH4AO
KyP+/sS1HbOaGabBxV/bAdOf4UtGOxb9YeMKgkn5g+D1PY8zRmIo2hHAR9FYixrxogi/08cV7eHX
fLIoHGyhDQRz9M6Dz10oluDkR5P+q63CZZbWtS5UM1FuzQPCkEQg0PdAAnlbpdHgM/VBgvOLrru+
FG7wgA9Tw+GPRvw1wJlOKzZ2WOYhVZQaYMTpGggyKCxSXFB+K2mrBQLLpnYuEUNUYzSkjbkOAUGE
A1+v8YhkSAkfWizH3gEz6nCyRnxIO05o+gDsdiaEAOBwKLZoGIe98j2R4+YO7uAVOZd20GWOCWKg
5deh2A/stUqAdy18ai8/Ro5tgV9ELuLKxDorHxmcIFW/7TA0xPGwVMe7k2iJJ2Ja0IdrDmlFT26S
WoaC6W4Lk/n0oUoHhvTwYqpwZ4WRp1LlBCZCjtfg7nRec3w0rqqVQGMMqtwY6y9tDZNrdgS1ZQY7
Agwt50aF5Fkbuczp7DvCrEs85SpjGJ2UYKW2vhVxt/C6HYcuxxmC+ugJMf18bi4iwOh70VSuABga
gmM6OjyaRqWTG9liFGIKGSjgltZuJV7ImX04WnCfCJv8QNcuwjbnENlu4jsQZORjDgiAn9v7zzW7
Yt0jFz52liWuXey0uqLj5wNOaLRNkjoyhldpmREW5YIe8G5iHUg6jgRqSFCLdX5W0/u4q2xagC3h
h2z3fv/oCGpyuWB0lKNc85i/pgqGcVoy1duvpqpzV7w4Gmvu9e083rDBZu3mKRQMCf62v8TLBXoS
YeTiENaDzdG1obzKY1Gx/DmI+v/tFMgAQ9Be0zb5jJdlt2v+RAehaCGIrb4BX8eTOL+zSAngJPrn
Z4WP5BFDyUJbfAVSOtpI9WfOQkppFOPUvTHXyJdR+idb9qjXwQNv4haLoIXI6V/wSAEJodbC9Xj0
sjd0qzXlgT9BBAxSeT5eBq9yk/b+OdxIDOBJI+IkUBb7SozoyO9siD+dclyiWo8iGNY84sIbXWkj
LV9Ur85STGxT0QxaukaF+LBBUYohs6vUYapPz8lIdIVILcX8+wHe/wBKiPDvk4QXT8WGcc2mCKQU
Ukw8FqP7uNt1CvjKt8Afd5dkP2yN7CEqBR5UY1TfZ+T0s1KOdc4x3oC6uVQGk1kq+MQRbIBbxuI4
upxy/f7ohSIk5VhEJE8i3GNz2JdZs8l3JuPbGUQbvw5LzoiHz1+rdtA4gZqhpwxe71XDOmN/s8aO
wgAhBfCuQyVuHu3SxPNvCPnpWKsQHjk0Rt1sTK0jcwgo7WzytLdgfN6iI2yGfLV8gnTsLGae9toO
et4xmxzULpWMEQeSqpAKMY+1bRH0mIE6zZGEdEiR6nrkncMmoNYTzBw+s85GsZgjemO87OXj4yhW
Tn836ejpYblItxk9y34t2NmfDBtw95484wADnqcZs/R0d8AyeCiwOXufEQGsGj1RIzrO1MmZ+M8v
O9c0B0b3Q52jDGUSn5WrzkXlnp/R1Tfd1flPMOxYF/a88rI2JNLcJfGTQC0AqsRI59ciIeOlufNk
myuicgfMUa2CA922rjjNWsvw8rsewqmzFgWqCFQjBGwawJHpuu3Mgj6asmzpSyMqoOhkOmGsjw9L
+yMXTXz4soPG9wtQp9kvJreZkjsQzam7VFDVH/+2PiFhFbIDmL47Fg9mZrtaJ4Gd1KU0sCudJ+AF
yhePHhamjANCrHHs2rsVaQC1BeVZhS1xQ+yfLAQbhFYNNxFNTv1LGOBw49AZPyGAEKX/b1D1M7uG
4OibXWqc+MaNi9mPYTt4PTiqDj3tmx4oIUzPhoNltKePsqLCPu0wz8zgLGCK8e8oNnt5fRqImVJB
c15f0bVzNu54Aqpoydj6lAb1wIWU++vO3sJ9T4o5umbAOSYCb3oZso1CQETKRlljddh7Q53QwwV3
ECbz8KXk7PQhI4nIGuxuJoaOPHH1vHU1K8y4YenArdKLnSiI0jkfk0dP/okSFKDLCF3dajen2FNv
XPa0QZhnRLPob/WLQociYt77PMKAAfAlBIj/HYQi1Rh+TP8mBz9eGp27WoKHqVzcaodnLHRILBf/
YzNucesT+RtABsAxw35oyj3Ysjt2yXnRpHqMPh1ofk1CYnJBdYCxDNN+JmwRJAr7uN0BEBqAF9xH
ELmQwwKaPLnYhDzT8SQev+6BoCQq/lLMaV+5AXJ7q81WxkaF51N+lwdTUSPBejZ+YON+yngNl3Qd
WRVHQEAQVsMZEN0d3encJtFk1kEAqS+xPxyKv1uGVpVja1lSh6MIZWWVmWEsEPQOYdTH//dcs8R4
meI+5EUL88hLzXL4SE4zp3WYOfQahL1NsJ+2hpkNJOzSiyBDOGfZe2i03hufjIO+0dOL7TcNI83p
LJ+/3fk0SdRWiT6Yo623/iBkmm9/TkPxQGNEw1RbgDWagonw5bEG2cy9Jg5hxRBzldUU3IW06OVp
h4oFPiNEmcngk3jUc5J1KfoCCU/F0xgdXtxJKujZijYZcFaqyyRyOfX8uk94CIaaHRQhMvghov+t
TzJbNi1WHr1P+J+FQjfJngQJWyff85UwGtSQtKF1OtKFwrp1auycHoepnqyilAOmYO8hsKQJnbav
83a+BCG4mGtVs+WEVTmzyAOiQ+mJXrimatrIp8SV2wEzTBeW1FAPCgD2INCT8u553JYXyGvc2Mb5
IWwp2Vktljwn61ucOkCa2fwtAWZLFDQ86jCIz9KIVSyRwM6huLH0etyHvM+m23Kapcgx9QG63dfp
j96EcuihsT8FLHfIWZXFk6f/NxviCcE4YVADWH7Mh1N5Qpp5v11dO6Brf2TojDfL9nAppX7OSxFl
U6Ju6F2JAUJ57P9xCP4+l8zF5KLe0HvH53g4qvXNou1mucpZz0vvORK36+q4YbDewOzc4s9G++AD
dUUYAGh6JOQT+2HfzOu8ugJq7v9ts5w0AaZRIbZQ+3vPoMQgaN2JJoVwZXHr67lp4Zvlc9HT54g0
2hTCzG7TXyby8PNTQng9GmEg49vtMCUc1+jUjvh5gbYj6caAHbzGMcDbzhXP3nQ90orPB6KhaFRl
bDO3Iv6ar47QuswTN+j7dJUallB0WAcBhPRTLsQYMZ76BYcfFypNWmKPnSBqbXapj3Qes94XWT5w
wqqoRjlOM/I1LYffaFjy+LM2EfhJL/f8AeO9K8Rp+mOSgMfcFTfyOwBPJWIgB3MBzAzF8j+Qh/2U
rvnLDpPPdXOFeTdXjwARRLCpfguhBXNNZ2zxZGHb3fh5PR8/xGrpcd/5z1fB6a8rY86iYzChi/Sp
KMWJqXAseq+NUHMmX1Wj08Xa9YMBQiHanJFByGoMA0MmT7zUiHiChFx3TF/2Ff2CUORo+MFVFLbb
xp/8L3Zwn4Kq8u6KFAtuE2f4wn1hInJDJJc5UkDgPMPo2ttscMHuGPZq7od4P8AJ6MIEijVUkL35
OTYMnRe8KkB14mAULcc/ln/4tnvWV0TbLLd5R3IMTwGDmIeg9ss9vZWotMZ71mmWjFhGfFb7krPZ
UG+gUdBAahILizjxQ/8qWNzfj1oROgNhk9R1uVLzYnpnaXOUPqODSJp6uGfWUvcC7R/htQZs62DF
/Qu97iNmZUrdaWuniT0HXpqwRoxIalCSMfAL8PDaC5pDpu8IKLj5vLDEAxXnmN++iUTfudj6O0Sp
VFs8rxSoP5Kj+N0/lY7vfPFab+TFU3qxoywUKyjr+70gZxfFarbpZ5pLNp/DVLvtbqn+O6eRTxWa
xl1gE9E3u2mfmbGKvgwGheHAJgQ6NIo8juMigpMLOpwHG0hxlpH+9fnA50lVDG/7uU/UM09b4lFj
G+RoyKOBizrU55BJpkbkP8Jz+Wzh2ki9rYKTBg5REv9Qy6AmN99bMYDF4MoC2gnSCbKodihug1qv
JaEPPVZp3mwef5A6MQ7hfOPBxCkhWsK//S7H/3eOCv1iIITV8njYYz8Xx6InoDyErOJ9q1yYEeSo
yPVDCcctIT6jXQQTIIh7FzsF4YunQaJ3KCkVtNzADd5PNJw2tRjrosXuZTTkx/U2laN7JZ7DlxHX
yy6+rL8oliaaS0m0LKfgvcsIY9CFWvVD5mFPqV1sQCG6z8dg5ix44euBssMyoUzA3HYV0v/UJYG0
Kdi1HMc/VkT7O8zgQUidxVyrAC1UPzgILhJsRq4KaUy40Wwr0RYZUPTYUDWnTPB6ftXkwtAtBq10
Mu+aSRzy+6yuycfQ7Du/l6EihkwBxWOaaTgvKDy14Diz0/SDaSqCtY0M5JFDuErRk0K+0m++Mztd
FJFKo9aiu72j/r0wQF1QcOTMmQTBnNR53Gb+U95hiOuW9fFGPZtZMscvSu/GMoi/ZZmwXv94qzYm
UVyN1MiSQ8c346ugQxCIsDidv9o32gEHGEyjShF5nVE+YHh6Pl2x1+sDFAixKiBUhja2/vl5SxXy
BOG72F1gBgfdG4TXIJHW/mjSrG7wrl8q7Lye3v3l8XzHTKHJXi+oSW0jgUlSfhlsQ5lxvs5vq3bt
LXNpWAAWzGblbfe4RlLvuBD1QA8H5z6Hb6c/oBwd7ep76deSq9WJVMy1jSrHlKoxgnQXvdItriEw
3mZAvSXiEFcvhCg62K9XbbEnfZqD3G/4kylX2YAtih0EbKcYZKoABoJMywUJ+KrAMQOCjPsU0O9P
RR9eu08KL5NJqvIeujlf8pz956k0AOw1ocFofHA96XvLMZnmxeYi3KZi04/EkeJhqwf+6doRpSmG
56IqJHHRWP1NYuOAjL5g093kFD86q9oWETVP1gwaoLZ/8/VvVNuN4hgAOKXRSjolZm4IokpaIiXJ
oTPdaKUvlDQG7DOVm4llMrqLx3KMylnsoZM6JVbJkZlbvY91qEMTsQK0gz6fjRDtWtO9Et/QQ2hQ
rQEeyVAjKB0f8Q33FdA7g2ZCvuMYNrYkDbsLSPpAGZ/8wkmhGHC/gVA7ef/Lo5wiTB+DUTgHUrEm
z7r0/u01cQH2b7c8c9pJJosd3oNPxZbo0fPLb+0zyBvJEZsPOeYdi/1vwdKVgYVizjSmRtWoULzU
LDdG//C/vqIshrQbC3/TrVQVMhmsmrf4VxsGmz13rQjiphYDk8Dy3xy6Uo/TwLbAeA+Fs8G5TnCW
FJklq1T5DlW+BfMrLcwsCUHThngmxP/P1h4WlJu4hzoP0ffBNvwQtD+RH3FcITjs5HsY/WcukcKU
6Y0bhTsb+uldgtTInRj68ZjnQxC3vSFglIkXbynGCiL5aocsxO2kcd9zjokKX7Anr776IP/g+OS8
zo/+y930At2nL7nwLqsFAnMApetI8DdVJrTYZBpjDL21ASIWK26mkNZWNAHyug9f8FCcyOqeFncy
kJmsznzD/1EB352Ln/IwKlk3rhSG/O8mUOtnkTE+fT2MMwFn7QlyP5Tfuo7mQ6kYfRrFxBzUp8i4
emBWvSo6fwXjjaztvD10ojEoVDuw/8no7KXqgHCJGnQxpORzTrk3SbjBaV0PmbshPy0uvraXHIfg
eW23K3zNOqXKzUFLBgc8YCwYoeHekd15jS7E+d4ITS8+6aepqLp1En/wSFLWse35rUzPa/fmYT6D
kkg64jxI2Zqej/MgKqUwuZD0VEyFdzri0gPgW17Tws+VHFFHU5/y4JeJuhXh5LWYr8Xj5O9TqAUX
eL78YSMxpexe54BoYUg2F6uoaBt8BTeXBiuPHrXnebvBtrZbqaDfoPrHkW2lZ0GWCxwDUg566ODe
v5hFFCyaVOMUlSSEDjZyy83WcIir6JrOGDxNnxzGwhqqlEmjuJsAGfPl/bhbRRKmVGFB83MrZht3
r661fvDDAG3S19p668PQ08fjX1y1SXEfEj+Tndo8ksbCRGKwJzkgQMMnentwzGdwib8hFj07mRBD
wefLIpHxPL4KELvh08Ak4n4PYMYGbnPUyUO119NHtE87t5GBYyEhklJhb77uCGkMk8Ez5Q5d+Xot
zXbZ6S3SqFYmTxy7V7NElkj3yB1db+am7J5xlXN12ahoLQq2v+ey3pRywjymA4cycyMuM0N0WXJf
kLL+0SIcDc7TVEb/+k036iAEieaTUf1qorcnbz2kkkZNQ73tZc4DRsD8cDE+FGuT5wCCIppiyLK7
2ZPT/4etmyTHxjm5cbMM50mibwjhOE4whSh8Mf5uwc4S4w0iIq4cpAyPbOp8WZHPf1ttPOy4vBCO
B2HUv6oqtR5kOIlQB40alp+3AaROeLh4MoSUm1zR/yKQGtDzCgPhfQPYKdBh+sJwYdVTRnuXaeuo
lX1jT69bzzFVCfRMpHhF44R8AissqMV881IrzvOA/lWAEGtwP1/fWBCbQSz73bLmY9geDmxUq6h0
w6hWFoL+CuS/AGspLAQetpqummObNRSnFit/ro+sfiTyEk+C6AMOFRdU9hmL78EfILxqahg3q6aQ
qBq3tAy8A4R1wSd0JREUrpFp1OVXA+H2gQ7tAvRscJEhlxOKDS5ubn+VYP7RtPijzs+yELTeEfZN
ImS70cdt9lUmDQyHkae/ktgMClON3dbfYtHdhLQIAEi5cVv8ySgZIsO7GZUNk9mhjMOabvWuH8cj
5KU1jBDBns9VXxV40doSOqG+AUGqBaTPkNL0BZcsIKXzajELpWzcDPptxrMKkydEjLB5G66UPitd
26/hGa5IRAnMi4ETzuBkOZ/sk2XH6GVOkByFd1TFf3wGS5TArfFiQhbOhTkbctYw0synZjIbY5Ag
+AIkl/rqVtF1GW8JXYwAocdSIcmQ6qpO2Vy0Ogga1dOWKxwaCXhjNZSB64OjHB5Wi8cSIdx5as8T
w5rky2Bxhr4K3Jcl3nSxQViP4OsRzZpnG7VEDg9jsgVZ93nBhMFAt5jxXQje3qBQKkutc/oc0koM
G9Mk166hRBU0RxAVE+pXb9oguY9+nONXD16YV10P8Si22eEDgA7YXb/GxF6hRnvg4kX/G33ibOnt
jCbbR0tdJzEDC9EfaRLeThk52pM0sK3tsXk4cD2E+MqqDxNdSTAjDN9NVIgJ90xHbgEw1DfsWB6U
ZjTYk5OhFJ1lcrWTM/s1/DAsgKoln2VEb3I2iRFhzZSAVJeKTUJxzPPi/gTMBYV0G9ou8jfeM8xG
H4z3YS2W9+xM2uvxYqe9Mrj9JEitpLf4US+yPRp/M/j9ovQ0qSz1vD/v713EgK01mz7jJ3cIDFFb
PUhZwl5RpBtm9ZTsTpMJwOfsK+csjMsJoXmv+1enLN+jZX95nS5OxJAvyT/5WXbxj6gfJtJ/fimu
RvIzozELYuESNITFehmQCQ7GR8NMW2pCYmAM90a6pvTi+2aLg2QtV2AE0i1tdp01WIp7CU4giS+d
RZV91dkk5Ey88pUMUSv5QW5zzLXjWD7aAlO6dQer+uUtort39ZLVZ1ru+xdpGopUG6ssnG97K2lM
nEIJ0QiuGuUs7P69nEJYIznzgt7qSYQkEdCCQCnW/a/j8vi9RdDtcN0d9wGgBmoUxmo34Q4QyO/7
oGDPc7dDaGnlzM6rC77uPaIr3B6byaVlokcrVOQSObGMCqi7lCeiFiGGvmYqiuQcUd2ikN41GkdC
Ax3NjDqSOZQEHaFd412SqPbU9OvsItEqxMsqjdF5a+HZbW5fH/GRIVokRh6GK0/N1sgl6X2jfIud
8yy5gkVJUr8lPD/MF+xmyZqOuD48AhvShorLDFJ3ZhyZglupSH9ioVbPlEEtFosSf32GmiHvtVWN
kmJuSGDIDKOf+Poqb9P4F8whu0ikngqIfiYCGk17f+bDgXxjbSk5WrInD8PpVuuFmVtWbzgarQrX
UY9kJVtbL37eFshaQyAkVka2XcYdiH+6FJk49Ho0PfyOEAhSK3ENPt9OdTc3O0KcB1EhKImeOw98
KljyKGimGHBzVuPoOO6HPjKX9k1SaDmdgVNAvQmGi3F2sgDR9rmY0Fsuk70TkTjT+tCmDR7/j9vZ
lg3nrEUw1WbYU+RsNVHhV9KF59GiGRt/+CanxrCRKgJKyVKF9CWvvkizMEITRkb+Zt3/IbecaZ/3
aeoW69bzjISUCiIYpMM2qdSpNdKGQo+rwt/nf4r1fYRJJdpXztFZEK22lGDY//0bJsSKv+PCE0aj
GQhmFed4glAYc68AGjc0XynKmnO72wWeJCLuf0hGLoXn33dLJCjGj0hxQePpc2UBPoT/WH332Rqo
hUn3RcNhSjk0V4YtemwA7/n8zcVKld2HExO2Zwpacg7gAnQBvdLrivoNSHW9gxqSdibRetYHu8r+
6U2Ss8dD6R1S/OaP4UwpiJjBL/Zjqiqx8qh1cBByLbXrnewXXiEM1mgAOwlcLVgr8M0v81lLf0Rf
aCl3c3itNtWkNs4MPuCOpTLxfBADvz2vCow9YXDZUsqjoR03SQp0PFK+6/Ma+xIJszj/HALEC+dN
PghviofDic4W/egYqwsB5G8NQQg+OkA61HYZMd7ui1cTq7lPP/qoYbBykAc8tpeRIjMDIgGN7EYf
ZZTMPugqquD88aTeDmmn3O8cMsbNvzZvj8UQZjSgcUaYoFxBqzPZy5wkfafvzfCzhGgzPO7blDl6
JQo/9g5QE0Tde9sp/Lv883Y7Gcxb1qrrywc8mttPaJr5FZBrn2qUrX/SAIvtH+dfOndOYEcDySN7
Ly0JBARzA8RatleagfJUKM1EDAohddI+MEmS2hA9juZumMSjkwv+bzcsUUper1M9X6zJl+UB8lkl
8cy9ER0cwAi4MTFKFMVw6xZMQfKBi5pVXZEPYyq8+9xT3BpQtdTPAHRaMMnn/Qr9/5Xo0KCQZ8Yk
H3baOWrY63A+Ebls4r48IlaYRFE8qna9gXHFXaaHqinaNN8fuPurHTeAdee/PvkNFHKAjYg6zQGP
8ptTfX6zcykjtY2BA8Rpb1kfChLP+TSvbf/QDNFUuat779WiCpW6hfrKseZz/ArLKFyqJr+8In8Q
yyHevMj3DLGJpNiaYV86z958EK9MiiSb3jT9rPNGxjeurfrzyaB8AIPxvdjuNqxsPxK7cPu+sYUj
TKSfi0I6cGpshumR7l57Mc52cJduZVNxoprLjF1vaLPO019ON7dEeYGNVKuNkQ4cFBxcQ+l4X8q6
Z3MSEvDz5VaknKTMToF3ZSs+aA0ILT1sCL1mkq1odjPPpdV5q5LipXFkUgYP6/Rxz9eaUBN7mQaH
rvrsb5aHV2YPQLEvaLbFNULtF1EIIWmuksXrOGPH7A/E28sZACeG0hxFRCU5wkkv+/AAfmqaWksF
ArxXUsc595wmTiXXQmTMmiwSraAAmqLAJ7cxikCZuFJE1q0//i1Hzw0fW+VWgqF40o82zhoSNFSQ
Rl2ccBgWZWIBDuAQlzSbVoLrvvKQt8jV0+QCzYHvdVa7GXVF7Oxq9F7lB0gc/O4HutGh2rB5o3uj
XwSFF4P1PUivhWjSOlDgbvuetoLyhephGVOwEIarNdSMABCRiBWvdi8KAonwFZq0eW4UkNA/S4qi
2je7a2icn1xzW00xVRzaZCX7DbM+7Olwz/hda/rqneSWw4rBX31llwNKG7zEhNy4RFgtcdRynCJg
TBVGLZGpt/WcmjlwzSftnv1OD8i1Zrp34+a9hL9fALilUjZug/o3yQ0lxHieqbxH2KGITSjhno/1
lT+8Bl2Yt32mAvMEJeFoSTRohlte4bIH1ifrcNkayhGilJ1mfI01BCbJR/c53iPQPY4tXut6n0bV
AidD0+hlxjQUr01Q9UIQeyRgxfMsSUbheNUkcT11funLXK6eotdT7N1CAurT01gppe1aium0ZLGS
Eb8g75Vc1GJTuX5dGFWdKI4SBYY1ms80+vdonRLlAM+STD/8DxbPU6QiZyu774na9shck8/bY4hk
XlmRZ8zX7CSi7EKA9ieheLJT40TyIdGhwzpO7hjLNlPJtRXuBQvypnIRsCbkrTyItrSjr7rYYo4l
rtSZiVAeonuUjjpVNbcBuGRfB8V6MS8Getc2gBZmd5S95+ZotnPefCvUG7PEcXOzIYTwd82ywWH9
LTRjMqPCMQ/T0t2qw1OAb7RZYiGEMPJmruyj+/Pc8Ix63hOfVKX2kCrcm7AfaleuH/eTQQB3hcgL
ZZihgGsdPjkNxmZkEkMZZ6kj9vNA+K9EjhHlthOcpd7jyatHvjteKaKLx2a7FkSvdXeOMtHXkLQ+
Ug3z6wLQiSvK/FQexkMfM4qFz3UYewbF10iw9TyjJYwW5pMAN/fvGqS+JWkRbuHHfgY/2vG37JBL
6iGJ4BMmysh9Wx4L0auZ5ygWK1ONRv2qERTCc+k8cgcRXZd1THwbdUjDwqUnZIvJrxnDHRxd3iWE
7ULO5EoOczwJa9hiRucMmFY12dNV9rx009yTgZ/IF3uZFtZGoPMivI9IeaadyjN7IADDyx9FVOFO
o7j0/ix2CZyu7WTEKHeYemVPUFdPGbzaDYKkcOXF6PqikK/Cv+TeI88u39Cf4+oa3DIaCjo2XlO1
GEyhaY//OroyTbdVELgYLpbs2q9z89TY1B3N9ceSkBRGUL04AMntTk0+wmrEyncrmbcUZZ5JSoTM
HEXaDPEJXWM76rg/uRGlAsUvW2Hhyfd8qM6896klbBcDl/ih53JP7pm1vlS5tdlxnb5y0iRECKfs
v+/gnrsk1ry0TdyGvQ4X4PHlmptMXX5d9ljcC7SvvRhr8oiBDvHX6YHWcMbZmiiG43DG3rYkEAAR
AwOor41puOez1d6GMpBWE1R93sHfk5t59qQasA2ERjvxBYjFgF7xW0UvkiZD/d6xs//2fUvkCqU+
uwPTw20UCwhtkSVtWbgyuW+FQoYlhMFhoBiCPU3gZ5h61Ijvh/KLbcQSa5dU38c7XqoPJCMsiznc
8j63KvaB8EbYrmL+DufUHPq+0FPj4kVyBKdShIKHXhboMeATECJLfEreBq/vRzYc/L8OFxgbmpEQ
bn2m4sSNjCOwle3CrNWhwJeQvgtkiRa+PMhKaa47D4qTWPejnYjn2uy3SIo/6Jqgh8lhFqOajGqo
gvsGYKqP27T556D/qyDdvlzcKEUwjdrbCodLGcAc93lXSXsa5FZlg9GVLuGhr8AdEnL/DHY00d19
b8+aw5iDBf46SOq7DrNp3L241/rJARaOmFvnDqNw9hgLckkc0fylXHlN68c7uKnTTYAmQGOehLJJ
vCjLTPp893AQSLgn4V/E9+9/AQLqmFxvWCZis/0e1PSs/pUDw7ZtvDhEVbonKiEz0nfvM1FTIlNZ
0voDUckFxybiXHQhlhb8TrIgAfZEGkMsJlZXZ///nbYFQiwWVgt0mwwanFDrgnDHoGVjzg0gS5Br
19DzRue3+H2+K/kY9c/btjNc5nK7E1oTLOZwuUC/dJaUc7mS+0KEYg5rrq1BF7B+M35sQ0rjjQht
55zlGintKe3Aw1QVs74+fBcofQg6Kcl6F3/sXQpOLuTp1BQjeAbWfJA8v3Wiu6zMhPUs/1T2wRda
qtZNNldaHmAvKJJX/uC3tpigcRYdg7On2TFNEa72BiYctobK8HxXZOLTcrxiwhNzryRCY4VtAzZB
E2qkEyoVkuFn8BtztxmSKIFQmY8Ua7b719+xEPVF3BMJHfMg5sLJLguER8Jp9YIQ0FyjbsmnLCgW
q3LGJAXXGvmmvQXsfRP6O1Hp21vccnZZP8FTmxvvCjrsY9/4nXQY4v6Hja5Fh+py90zXRCKRCKTU
BUV3j4V6q9ZqXyW24sQ7kmXGwzTcf5SnNYDflQnf0nlPLw9wRGT/vz4hlWY/xWEsZXIESumMgb4L
KXkIaLVx9ysw6c5h5VKqW+wQx9jRlbxEf+uJFJQ4JvfkMgW8FlEYZWvgKXNObys+71d/4wUhAAil
OZiS6MgFEcgMSCzcrYWmSxgYVR0n0OaeFLhKB/IZ1GHmpKmeY9xaCqo16ao4L27rWsQvE/aPTYtj
kS66pk06qAInBNgVp59mU28sg5mi9Hb82mTL48g2lKBwjDCGuFXLLYKerSkz2PUAfgh9DYdron9W
uXeKFvplh7VwfmRIFsGExUREzD+0FMpWzkevNcTzzOZ3sH39wcIoMuODDuS9qFhH9ZGwBNZ12PPH
MSUSZwdKwpC37Xa91Ij/Gj61yOWlDN8BR6BknOf8Yq5e0rfvhB5Wuatc4TjIF5CKKTlc0qMgCGmN
ElyrWzDZPRuQ9zbOOlHtu3Sn43cKI1GivMfKPquCmXbNupTHkfS0A3ke8/3DyHEkvitNAy/T+DdN
4qvZIe9KRbaGioZkZaX/SmR+pLhQi8A3o5oyFR3QQNQdU7OyVR4RedVLsBpc7Yx7IFrsg4yOqvha
n92fAwEij4dCc3gI0q+a6GIYZlJ7QGyNJFdQiCZLCKHr/SVFQ2azuV+o9qqEijD2n3qFmFtrqD2f
5Px+txQKRYOctvKoijrcew/zMpTKu8FGVk4Nsjzok9txRWcL0G94MrlnrCzF69Vo7zaxpAUT78i3
F2XdERyhrvL6V0xJ+DQUKRGwKroBOdAC2W6fGn4da1ye+mND1kY0hkkvbwv/akNUBWkNILdL99q4
TCESHLDDC/osudDBaLyd1K+boMCF3F+iz7ko5iLk7QsnXWQ8TuQj4OpGnW0y8ysPcJcBUFtwep+s
zemBgjjZQD18ePu2BGFNnOASbgFnWu8cCdHT+SiteDU79wbEym6MnbGch5mZhIiDAB7RA7RSDwhE
c44fufsdEHUtfIHekoV6HgACc21jiCsXQXVTzV0bjgneU9Bz1pnZkPr4+IDVhRQGuboJCgMBhQ5l
PrPI8sFllV6hveVp9mIHihrxf+tpjGMr3iBV3CC/dtJ25ywABz/L6QE18cKPh+Upy0lDAytIxREF
KFFS6yF/rUFxWM1T9v6M334bVZs4/YJI+2nmtOTVd1CI6tVn1CHq7llyzRYPHDr4CCASGcClEDPG
P+WKW7PrLMEP4CXg5LEFt9nZ8A0hsIvlPJ301Ui5+YLnlsl0vTwMeT4PspyudtQT4HAJ8TKPxQkI
kZK8mmPxBee+GG2OR196qJt0TgOUesZlJst2HQUlFc8Ljs8WfMiB/VJlP99m8qKEzznPB8whsOV5
GaDVnO1IFzrx8xM8OYTj2OHRNTrN3hmXneFNvMolehvKGs5pkdo6oWrlsubC5mXSbwKU5g891co1
24KfeG3JXX/MInN0W2F8GE/GxDGkZE3cBVYUVl81B4c8tIJu3+I5PTAHEQBhicHOl/UKL2EMn+bu
sAYcd+TX/U8Xstr+Uo9VGWPz4A8ZJ92vceLfnGZmNjjvmjI/kw8RtPOuxEdTHWFDZbc6fz38fj8t
JXhywOl5eElMSYBrbRsY6q9wTsbplcryvKFAunnWM5p1qKLrmDy1ZFiPDhK/ZppyJFX3ea/DNU/f
Mij8hi6pgbSUObVwWdXfTojwXViRVuPVhC3RmhaYdm9VU1okGL2KqN0gsrUw/L5GiyxUozarFmic
Czqho9roxpZzZyHWd7A813OiCkorXRDRWO65iW7EmX5IB+dFQ2W4DTeXJLWFKU8Gs9lA9n8o3/GI
aeT8xvkYw4datDKibsg+AK2RJYS0PnlRgsAuJybYNflLc14kBmAIKL57VvRArkFgdyYRUIl2/jVB
FXGfDsqiEIEa0/cUrHSKQE5PbsJJoAhFIm9Pr0SFYWZuvaYZ/1XNQD5G4d9YInOfQ0uXrEqtcYQz
t5UVyB6zt1JCJ05q2GxAjV3w9V1H+UBs5+uiSI2JhGfFtLbiqPsMjzrLX8ab+rxICqFHWP+aKfoM
BN//Kbi+gfX6geXKBT/iTYFLWH0hYfYY/im3lsPD/RqCSr2rC93RLe3tFCot+Dj/QOsqkPOPi8mJ
alq52dMLdl5S5r6EoIe5pQ7MwHlLqxhrdgL/kZPYmx9ofBYgRf/snDJm4tytN2g28475EsZl6ful
H2VVaJBz8f2hjsrGxushUmVU0YNPRsFG14JO9MTsxP/IttDnoGd8hgB6QjRMheAHEZ8IRGfTF300
gXJJpvFo/5bJyFo9wYGNKe9aYF6nDhf5Y/mZNImI0TBtCz1tCjjSZ0v/pxQ37l+DXukileBjkwF+
Gpq/Ph81vMull2pYsBc47kRnOfcYVPTqcPs/WbYsZu5lQm5/IqmKZAB8LQenP8KXTYoB3iIenRi0
zIRi4/Ew8ifjNvX2W4C3yf1qQes/YPrg9JFzLqtxHHGk2NYSHMIBwqYL+6s489MJGd2aUisjphYU
3aGCyZG3fGr2AqbsHYPpup5WHu4qNAS4TjgpEJsSxa5hxdedPKI+QkjWjWvNLYZAh25INs0GwSz/
rbNSrtQTUmxUnjrMO/NflW8dhKU9YYJHvQPsjXWPJpGaSdy2yIiSS/IUNf+6BlQKmF6ZECxT7K/Q
4VSJBQcJyiOZqb74M6ftOmIGiBZZQQG340x8Tp/hczzjHMBwaMh8JRaRhU+p5De6NcLXaJj6Q4sJ
sb2VglmgzBVI8Lg8gcD92edC7TtowD+jd8inU8OCWVtpnKLjRQqi4pJuB9GclEJI/D0sXif5e8/m
yfvG0zTZEmKNrMHg/+aJ++ejvASQcqnA1WF/Ko/KFMwOpo703ggoE+Tk75Du1EXJ3o3GkjHnQj5Z
cPVuiAgEI6EhU30yyXQZ8Mg2oRnf8kltRPnp+rmibKQwu7b2ah5RiqI7X9wV2mGa95O20VLyINop
SZTCVAvX637VbVdwo6kSfWpkw1DpasVV0CXMQd7ln9+fQd5pqN83Oa0z+/PjO6eBXoHQscBQR+0z
i7IC14BDxdKpSaDOuGgnLwjlbY9owSNspxRo+sFkfkdbcr6XnRJrjPxTQVC1ChAkezW7JWpAM9XS
Wrtsa8GAZWv2Lrj6QQWsHz+T0NOVAA5lVn0MHsiaCBgKnGvC9xf2TdqRmf7rPLlkBzLg89uey2qV
Xa7dOK1IZAAnew2Xhin/oKiUB0pWCaN131K5n+7NX2qj+DFrRu6GtpBxkPco/G7i1ACGtvv8g4A2
TmgpLyQq7BM/KXx0NvSrlCFWj4vK0xpjRlLYjGqNL91womXMZZA/sorEnE44Hqpf17RYk8uCZ+3j
IcpGdxZPTVUJcbwEfvSMOoi93S8WY+PkuCD5hMwfZPKgZp4s3x0Pz4/MHTMxWUeJeOthxijeiV+N
wHQIqlNQwwa3uhb7wvPIzdPLTZGDTqwzKeDyhfKVukDCfQUKi5SovsXh5+3rHP/ei2XIQs8ri3lh
T8KurquDExRl3bkmAj62R9iXjGcD63PWbanri4SLXKMk2pUOtXXtLur+fKw4raYu2+EdJgZu09v1
2zv0NK9fufDe21ji+gG7dX9FtE+64wViALthy3OF9MCZzVLaSBvxyXRZ52Frx/v5jNxjCbZRlxnh
iOfMZsRDwImZaoJukmS+Wwc88jDxDQgv6Nq1I3rdRx9WQtRK3SavDTj+x9ghUV5WJGv95YpA5tPI
JyjNpFHxJbyNr6gBRReIJMJbOoUMIKDkDfseyzhx9a8fxkRMulrMsoZ2vKP8c45hAXEFy58qU08s
BPnlP6z7TWbo2g7Hx/IDv2q0Hn2zDy6F7pEnXuCkNSP1YVT+UAyYpU2FMI6HxbCpCXx4w1CipPUZ
EcFHNc6umHHwFrtkjiqNiI5R4df3oK7AbRoKdUwCK5tpfUUrRxZN3axMGv/aZVvVx8mZ2dT+MoWH
jmZkwe1o4dSzew3oFPhH2FOmrth3johmAU1zQWTZd4F4bN3dTv9C3vAbSi2tvThzLLnHAhub1+TJ
3ulRgzL1PWtoW7ULgoNHMwps6LLFkYLIEBVKDev23QtLemmlva2YluGATe6XuWmlgPuWwgZn5SWk
cKTSuvTntxKJf+Ru/77jTIiglx/Uf2Yr50mzkVW0s/X2AbjdL3QrkIfutbWKqyigEMF0Kk6GYqxV
954+AsD3wO6qGprEK8J4MuR0fUrvoR4zx1po0TKUz3CGcNTFTrLbCHM+eXhVJiy3LpwXNN7Id2n4
MPm1pziozvbMEIVKN2HKqwZczz5+svlV7Co+maN2lSr2j76/Pne3E6YYWBtm8vtr47IVwsOD/WP8
NZpScHWkZ4A+oYhPDsF7IjyBzW4bWR5F1qCaO0CGwDW/Fb9a6k4RNwh73PGmBp8aneYbNYExNfUb
5UsbJZ3nX2hSkXkX9X+oEBnapaBe3jkvNVIHlkCuI46P+tSAcbP+mPhY9dDNkNfSwUoOMrl9z35E
QmdGWU0ds850Szz3tZik6jOrTwpbI6xSLHbNbCGLqQAJjICqOgOFSos2m6TurIyz3FYEIzOUL1p7
9LveoDugDHxxYkxvkeIS8w9VYmdATeBuwz4zUxfFgWNpBJqzOA275qAITurQj5i3THgZqjGge/vY
cYrDGkopkEQnmeKr3ndoyEFMckwje5qRDTwp5Z3+/SDOr8YvIpZPtFLFDPmLmx2VNbhkWrvIs3it
bHz9sUHuVvKkhKtcxYWOeijmV7PtIMzb/+pYE1+z6xSjekH26v1BbQI3d2d42tip5ntXCAtXyZER
E3pfOobjC8BTp6TyfSuhv81K1MU4TZz3ab1Qb7Ed/ItXFnN3+IJtmpv0O32OG9N7gwBWqf0Xba3N
9TFP2I7MzyaCnF+cKHB7xNgOXKgJmGndJc3cpXhYVOZlSnbK0CahsbpmZdyGf6fFaT7EAOiZH0ek
DP9/0EEnZsfregRy6I1U4xJR+Ew3wb7AZGal2Dilt1yPeLcDw033ZRhh5gX9gtLWGUKOhNGqHpFa
+o7l3P3gjd3U40ySekNO5QmSFQum4jPeEgwHNzBpuZWxkTBJUeuqeTEupAc0PiT0Pn+SIok3441u
9cIuq+KFW5zb/5jHv4KW8cw8dZJpIdJg8kGO7nwdkXWOkDli2+qvHGqOX5gWn7VvL1TX3U/ObFf+
+lcNy8REfQwxaNvhACp50T+Te2Cp2Ir+sGuPhqjE63CmVrmKPBUST1U/SY4JbH/V6562d7myIGQ1
/j9A8vgi3pofgCm5X4A9UmVCHbeQR8xvh8sgk6mkXrB0sTpatkn9/Gw54a7BgxwXOG1keLybM2FM
s0fUcR9Db8IP8+mNKy23BVx271nO6iDe40c45SZ9bh9cf5k/xW948vGtBOI1NR4qPzRb107DKTgI
zjNJjQFJfTjOCETjtSY8wORP1kgF5GfdmYV1GuBSnlvCsA9QxMWLYHaXEUQDeSNloigRedqK5xhf
mMreH8gIDWA0v621nfT7zWdS+zU0iO+75mptec08oH7KOTNNE63Awv3Ea3VAGWVFVouLSeD1f4DR
WJkqnf7gGyLMlfgEognPYmC25LelzE1csJ20s7unmd0+KUdVXnRcJFZGra3QLC9EUygOBDOt9Ro5
TBWBNAgyWuL8uZxxiwawUG9airgQOlmX1YcIBJtd48BkhZ0VudxO5gpB3chL1Wx9CKJrKKZp2mtm
fH4GjkikZTZNBE2b/VsjPMdk4llN1Ip3HmtL67EjgpcNd32tr+E7khhIJSauqlvq1ttrWc8yN+g7
qFOtWQJy7s5pozrxtxJ1JnDFy7W6DpN6k71rXznC7V5MKqYBQ/aDxKxmMfao0sIRpe78d9veX4oJ
DqtPXmRPFK1p/4EjaDtYvPACKRUKiG+7/QAzs8moFxyuro5FoA5wwg4bf2qNuu6+qSVgWWCIpP2/
twnylt/CQXLrys9DJkjdOn9e4ei+KhCos1K0OqVNQp3P+Jab+rHMIYDtfpUfup0cF/eSqJpLgwNj
MIb/NmmjfdVk1amA4wtQ8M4gQP4GCB5RDbXn3CcjvbwgZZ4+Xhnazj4+70NxudIgSd2YLzEenT3S
vL28A3S0Sg5XplevX6B8PKrhdh6oP6eO1HRVWGEthBihLrfRQisWCMVMTdTZMuUEp2g6wnCly6uw
P/RKiaej3w6B6NMJ8dgNgdVlhnVADyuY7/EFQHACYAa2yUtBkNeDUx65t3I4R0m3WZC+NFr2eifn
NuKro8gycetHLJmXd6Zp5pSq4h45TdhSVWHLHj4nNYKUvHkzyHp2HFaJS9LhJGeNIhZuQX2wpfZy
q00U9ESEXr7H30TCDTBkqYhBbmkZGcAvQP4e1StoOQPdU9wLfXGizIM8LSL07BysHiGxPP0BBVsu
ISYq/NDv7tEgmNklhM7cf/8D9UrVIce9ILjNadgohLR5iEwNdZHICrmezbrZI3b4zgyYLDXVzheC
9E1M8EpYJwgMJnDaKClcm6NjUTs26BxtsObCJADWIUreeHTpm9ErZD4SRVPnBEmHL6Mpycn06vJw
icrrzOqxyW9Eehgw/7F5Uob04se8wRrWCvuWSauWua+uISIfXQhV3DzuLQnbz6lKPZ2PWl9nSkZe
K7/ZSvZBi+Cd5IMc+u3hEuYpeWh/HTJkVTYlCCMs6bvDmMyMIRr6IUBycQnZjhf0Ow3GQuf3wuyh
OrU/2HKtHsZpI0FvxZzkALx80bOcqarKFQppu3b9bpDR2OeczoyIV7dIPVDjUyjQD3FqoLBbnY59
5Qtogg1zitmmunIErdi1WbE5wNOqVl3mgMkH25/eQetZvHY2Q9WzlJJKzZm8kvvvTAPIUK+XwoBB
xqApVMcsk108ZCJBUniKK0NN4TF7Phpz+a2/F1OrwOQcB/Hnkdd373HK8zbNpLLAhRJdbcnRvYSE
7uK2NZov7QkD5oqFUg8nUnqti09eAyVNcdFYyCRfl3nNO1PSrjxCG6/DwrY6jyEkRrizgyOuXLj8
+gyS4xSyyJc41jAv6WBmiEcFdYvFubN886zTb73YC/kp5BBIy7DxqD/fNcO2pTTi+gf63uIFjKnd
M8y69EVG0EQmR9bOqn94w0yx7K0pAyAhXE9beaZuAEtJGusrvpPTJ46Mvm8XXtaGZ9ssPkGfGmZH
CMjx0KD9lj/5janmQmrrfqMFWxJXY/Y5hG+f4lVntcSQhx/Nfx9fVJ5/e5PJBcd5Y1SqvvbSG+KB
J347KZUh+BNhn+bxaSDLj+X8nXDEFrUTTmNJlc5CgP1IzhuWdardC44IhYe0NcIFdkHxI+XQfWHT
tP1LUBDcodUhWSoflAAiq3ZFZZc/hPMXnLv79bCbC0dERQwg2JNNEzvz+aeu9IrfTrmRVEZmz4ON
0n7VtpZIuD1nBqaTZ6FP2np+x1mmFLsR+xjyybqXbOi31l+dZHeErVWVxAiW6P7yVKNEKJDE9Ahr
9aomeLP9wDso6E2xBwUJ/BQbwzjzIEF0+/HFmW/rCgGpRmXE5JYoRUAT8FSGRlwQ6jd4CNh4HYcM
GR85cEW30uOB8UWhghNmX/omLEdRQna37/jzMobBoSILUMdcQOtzvw0Wwxqql4V6LiSlAkJnCsaH
1aOm8Xvij3j1Sz68qQY+ycej4QGu3LynxYGzsfXGKe/EO+FilqgRrntOc+iUn3pQiRo9itMU2v1g
T8hAJkSlujBWD6HsFo/FbyK3EUPXzJQcbNOUeiAKXMRqMpr+Gf1tv0FqBwHsYgG6Nm57rkWGdre0
uWrz238RcUBWtQsLnFP1bg/7kxyYQoAtjW7PL2XJQZZHLh+1+XuTnFcCPS3vElsrNElyzKyy3w2H
QYHW/0PiDXRSXIhIttYf/Lsgstsu8KkvanhlsKWDiFxiPj8qV0k9gPQPOzfldCH0zQM0SlT9/sbN
i17F5DJjoG3OV58kLHjVMtoZfaF8eNATyJ36erKwBO26eRl/g9g1xeKYjGR7Ok/BGVt/vnUSU794
tqRRaBupSTv/Vkj6Oz0ptzNb1asfqJ9hGiB0XGDKJFjp2E3yBT4yAwramwUhDeQqluHSicWVeKqA
WSIsTCksyTMlj6Ef6nMyE0NeASdd0op0FUlH6NNM1KJD8URvIsuNHiMahV9aIO8UgsejoSry2+S1
z7cqRuv02Tn9Mpn8QapE8RlH856QUHS6QKcpcHlQE9UvWOngMnsQrmeOkEvUgNcFioXlb/VluCbB
OiZfqUZoUy1UHQ2pyNuQXkmAI2DZh6H3J4uQRGznekeYS3ZbO8TjH2wvsy1/af5vRcaP9Xn6C2wF
BU1gnP07anPa2Soj0lvH8t+K+dk3E4KK5PMU/jzGHJyLdTjJOUoAI/xONeQh6xMp0ZDLX3x8SMEP
PChUqSx2UBHIeaU6eWymaC3G8MFRIYzJpMOwecTvYzp8E/OXyQlTeR/xtq13mbsbNBgNm/80MC2Y
NsDRdCZYBik6hmFJ33fS0JNZaTa/IrieTMl2djfUXL4KXe9YIt65fuj3RCAvvOlPAQLs6EZK3z3i
zvqAyKcSf0SY/Fy90XMrCssfaH5ubUo8EfSMpS98nOxqH+v5kQZBs8mUxmJ3WuYkMux/CLK/ExVz
r6PbM/jyjmt4SSj2Z7SQafdHeeNcOhBY+AY7T/Xj/KMaYZU3P4tA/DJ3y4Jo+DyWSf8/hb92Tam+
E7lGQCvc+hXwQqBCF04yCZslCZJCbkGmNvs7zxMcHq5w7CaAguCxPa1a6XCX0y2tEQzggVVtPjTg
GuY3JU5NKtXlUNeSD0K0d0+vGia0X/LforPPx99QGE5BTKUvlsY03pCVLntnQvk2HsIVCeaqvBvA
xwP6gq1DAxy27EuepWM1YLoHZH/fxSeQuGi5km8C/gYEANlpZInPzOC6NuPqmBvPggS3A/bsknAp
Og+THX+IBKypYksIesKga/YrpwsgQ8hvcMzgtAFiIYpQEpeoLqRpxKDqvii+gvoQupC2o2/hLCRc
Zp6uVlmO8bqkVaPPSBlb7TU00Ew+JXoNt1aJWhvr7lETMQnIV6bV+wgj+3EHNWy65VZzQqHEh2UQ
jw32p6q29VKBjDTF6pN5T4n1ZyBbZX3uRYFSk2RMgTmZ9B6zWAE9ILlYRLwlqKoW9+dzCgm9gDQn
idLqSnJ8dcGn0RaJuv7xwwn9SgOEmUGUroXhmkLIjsFPS3i4Xs512G/f30ZgIUjyb6EfV5mmFTiX
+yZ5i5W7M+0khmIcScElhzYkZehS7j9gq6sk8nd2BbEaoutoI9unynOTqaqViDCvcVMxlUA397WT
Uph+LgNXgildFhhnQd391QPW2P5jNXVCIPQ6QZk4fUds8CCMwcC/e7A8urGAhAcVLy6UmbGl1/GV
klLvXbYLQfasA29l9ogplxk6WTebVpxmAkQHAoCqIjw5vor9r6NGR/ujXdY9Mv5w/cMWkN+Lh52O
tuzXJArQ1u3y1WpIrQehzjWz5SEvikhIpeFSb4Mhz7zboJQOkjCTl9DpuAF7Z3glAdfmQ/eV3tF2
8lSSlUjMwwNHpVzgpNxVpyulmVbyWpuc3DK9qmQJzszkLs4u8/zELQWJVTu5b5OFmaFq2Fo7mOhl
UMnZU08hhWDJCra5pft5DIzZqYYk3ie83SO2Y0UXmxYto/2G1yoT+9R2ydDRkgxchKL1GyiFMUDe
w6ZcuX/yV2tnq0CrMrKgtvPdBQoMf408R+QvL2jy5nq8HAM1MdFJUNtbeS4Bv9thEefQqyPSBNah
HqU4DWy8+ZV8MgYK9XCjbt1Hbc2Pxig1AdlvUuv/tzQ1Cnmrvz68LYzcCPlQk9M1TI23Q6OF6gk/
q3aYxr5qmSN3HBg9q+hUTyXGtgz3UyLrdlzqIXsZ0f9FePjdcYgoDr5I/ljIzpUl8krwQ0P82Bdy
OVEexeM3LKdOw4Q9MSYWn0+GWZOKu4pznP3CfUwrP657ZokujNdjBfkPcae9ooER5zBXlFRq0PQR
aYhPOPLH+6e+C93+45EzFvA14rmjmh9h/0W2gazODw0hpDoWtI1vhv48EF5giD4d41rggIso4dw9
9mgpbi9Dg1iX6TmqHZWa1ejBAhhZ5ZOTourFOySD+p8gobiB4q9rOE4lKlqUKTx3vvU4mhrwHNEd
WyiEU5r+KUwUpxEADH+Xg27JRyijrSs53qbvkoIR6g/zJQippjX6p6UDsNOO/1nJFxuko6NIet08
J8rAILB5OSfQJ54ffMBHGiznltZoXSBNlQXAhX74WbUJjGbRvm5ynw/i08BqjBVpN1fZRyIoQIQ7
yLO9yM3Xb/PWpet9rgj4kBpH7KKUsvUKhohGuIs0OA0TO2o46SxPzg9op3UbpiajQ6J/1fMgqWun
bzuchDFfut6dOwh5G1ya9M6BTf20YYXw2CHb+DoFQmAGA3z0Z3dUBw9jpdbr6uA6LmYZovFfA7Ck
WzNm8X3HM5FywCATP4yq1Hzk2kqC3fiGYKlUBIF9mMgsHGSahFQaIsckZxkP5OjXrrXjs75twGcQ
RTsLmn/heSpoilfbmYQiWAapDK3UPt6I0bXOD3M7FHGgbIkkrytH6HJ/lCgCCGltvMjPXEfSTjCs
F5lkYjVmziCoUkBrImbNmjamXZQWIG77ocqXBL5M7X6QvwGV/snjNFUPrlT8XC5X8K2mvCRR3CrG
M1ctDBMmNry7FgXBovdqRS4CsVYZ9DVJv62EfyYeJLYmhCujYGBCopeW9P8ZzTOX5HLUGqhd64YE
c8uAFXgHIPX2cO4TTYw73gDeNiDsKq+BuLD3FQOL6jdMUtKz7WX0Mx6izPhcSCMH+D/IF0MsOFVT
f6kTEd5KunWt2CeayM3Nfx0DDYyQULMzNiGF98khjezmQBdPiDSIBFg0fVQvf63Cng4TVbblMO/L
QTdGrdflrS5JSVBC8APW25KybQtnKhytMky1vCWI7OFOSj5k0G7A8js/CxWd0kJQjq0RHeaDvafZ
x0xERBjLEe5VzWo6CAp1TPuUP/JONhdaprXenzS/Adx573pZSjiCtreshyFySPPoCIaGjMU9jHRo
aBL79AE3OskhGkZlZvHTv7pNffEdEyxIvkJFtfS6PixwK6yXKvUhwYFywbJZPWoGWzCUjli5LLHp
VZG6wminlb9OsWmeo94pdvdjbvWR+EY3PI3YII4slrCDG+i6D0F/6IFx3x3fxHnpo2z8MhDhXAlk
MZUNiRVTjfpbQW55GWrhhyExHXLGq7lqHUjrHoImJWVbXjwYlKbcBlXu2XbIo1yyhq4zSkY8TrNV
+LPENu6ti+X6Fthf9rZoWjREfZFr3xqei1O3XjEEdi9cLf/54ubHEmk+Cpa7UdhN/APTTAtafcrW
ZyxdsNCg4I9Aooz/ME1lgk5tDX3HkM+Ch0Gx6n6zmH1jS2gzbjPrCptfoXItY69Wpw/SdPeZlZUv
itZ+OGSs14fnDaGkgfuPI8PVLoZa1T9/T6EWOhhKFytEDTFIjRInxEhP+0dCpiwlRINOoyXiwTf9
vvP5Mi1hI9Q0kOMusTa23NyjS0xE2QBKV8CJhpEu3VS+UGc254j9X8JDNsYWbDgiDYXey6M0KRVj
9Nvm0O3LvC7Poi+juCI9gp+xEx5wrnSuxTU3/MCY6Lk2ipI4VjI6ZeOD9Cw9JgV/RgHjTrVUF5Ji
33JsTy1cSLDRFv00W170nW0gWJjXBmCEeJl4RvFyAWDZVbNGGvOwQ8cuFJNUUgvXhez8kZAMnMyq
albmsqDXz3qC4+pkucEFTYjJ3+liy2hJ0KOnBtDUN6j+JMtM1BoU8pb8wbTjx2gXO6Qbkk+tOW/+
Dx5GVL2tSDzR23l9Q2VMrQje40Tj/exlIpRNVKnldGsEOcAWCosLCSwzcVHCJ4snV7EInc+gNgWQ
kU1OMimiwXc7p644X/rtDsic3dqbuLpwC7Ndc1UnpIK0ZyFbsMrwxUSEc3A3ILu2+P6F30rgDKpq
1iwNN/Mq+WBAjMvN1EmCVswvDC6tSEvqIAmu9C7FPhzKHtpzSPi9ioJM8AjjPQ4hf7teJGLN0NEl
yoj7VqQ+tHknDWarlXncYoMVocSidOBpz/+AVPhmn94pxeGWK52/wsnsiz53fiIzDZdcqCXsQVCE
6S48zFIF/vMDA09H6t6l1mWOoSaxuc8xcbwxYQAUil/1R3qi73eNU626SHRpP78fmEc5m75PUMCT
PT+nRS3+cQkAK2+vGX8FmjvKefNjCfkiPXV/P/QQ3qwHwqWheCVvvGpmyoJlani5ivcikEgy8nXT
k1dfkFYBp/HUEJ7t8LcmQRBljjHaEWZnwuMNHGt5FC8qxqLLq2TCi0YA/M9bAbdWb1gfYUnLpWkl
er7r2zVpIcm6sOphWrGsLPiP/V5kkJmW0pVeChTqugHze3OI9xasizOJ3wZLmDXIBLVK8tMxKm34
WgBdyj4nwW9MzcZg7stfrN+Jw+xy/bVYa8Qw7hnAfKphF0Ox5B4mpia88OdLqcPvts6znTiMxLGj
gwNsxMj1prjN/sAIBedqQ0wctetdQoMBY9FuyCHxTyM+nSDPsEJIzjZjHjc3lSK4qlKByjln1uiX
K6NMrAI6q2dDlNoBiMTgc1UKBtX7WSKRsF5zCy/d8UgspGVjHTHzdr5DfW1XGfgi6rDGwGGMh1jV
4XjzxfBWztIX4Gj79kaDNEXIRwQ0S/339ffq8pcG7V1Lz9Zo9T/BxHsUVFHaRZtHn3K9GwoFVzpC
x9VpIjJAak19BNeeRpn5LE4fYKgE/qjy8ssMPeSRO6hsTarmk4bpqBqSciD6QzkWskhdwIDoG2fT
ffOm13g+BZt3vb8Wu4bjvrgfUzLaXh+NDjNEuEhIblQKRyqkl3o/m/3wVOQAin94EheybdjoSYYX
vGkQMjNTnr5+lEjhz/zC17jonysisjEIasZczNcBL3w4i5ZlMETt3/G/v8dvVqbdJ2Mu2jw83rLC
WaZE8SYwrbiaXcGNIBY+Rtv4jUfz1NCRIj4MqDx/t/Itu+sq1P/Syo/9YdnNnqlLTfjYeSbXIh5l
A1C6gEhOaHkTEBwxEl77suEqc6JUmeKKvorVgg0uxQ3lJvTSrrc8nNDAeK1ItwofbTnf7QgyCop4
mBfk+fKiq1g44YKUCYTzhPbdhjz4a+gAir0sG5NIE+A86h7d4YUdUgnCh/PUAeMiQVOlYDWSiyGL
UTm/bNiclWYjXG6h5QQXYzWzZPfqN3flucyYJ2W1KKYq/7WGOvCnjxwvzQhWM/YaSGdEJpTd+Okv
jS8C+sR78R5DXNF5QpHYR43bFGYvWqdrCEw8T540SWev+Q6ZG/Ocl189qyRqFRtz83t0RfIc6eB1
N0QuJTNUZIkttyTT7RyFePdvENP9s4ouFN2rBoMjqFPw7FM/ozNpzpdLe+BnoxeNI3VXxFubAbQF
uzuvupxM1RJDkSS1gUJEZx1eAyxcR1+SXgCYniKTdE6L9zMkHTxofAEyatmACsTvJ91HX6/io4/O
IpRzlahTLIo3wmFaTSfFH5P3Q/nyEo1QY/+Q/4WalL/xXepUZLU5x6E3trgj7CHybPNjHeSTfsQ9
Xpo5F43RNkmLW8pL6T0tM1KX5UIB3SCzYES3zosYNJ6q35H+EW6Nq7mesQZWkcoXN0Egq6n96cpn
+wx0NTe2YzPwHWzoOj8BpxRFFMZy1GqZGZHa/wttjFgbpQLoWVVE68o50T/N8hJTtOSABEIpTiox
cjgN3O7xQlhOlMRdDIPrJ7g1adjK6Q9PjdtfKOcO/sW/CoYg0N2PTMpB89p1662V7ShnFnKIpDP2
TJLHMR5tG7adseTDra9zgltYCGDv34YPuQjHHDDiXEju82nG3ku1tVY2f1T36G/MaCrTaZhgsrYz
SLlIX/4hm1DTYseOuzTHP7DEqxdql+joZYVS1Ljf73gdV1FO6ElEFGPNyyoYPm4wNRite1zqI6bH
goSK5OAihXnhmSfVg5UngDaCVqQOlTu1OpDT5gSaAoRKnUeIw85W9zAwMZDPrvUnZi9q0UFF5Y45
TDlOaRHpR0mJQgAS6/XCVdTuVcqykbV/KNOGYw1bqw0mNRZacS9WQ9uUTCiJyzd4X3xIWFhsdYRL
chIQK8BUosbPzOFKTBLvOSDR3DBsRPQ98qf5MhvaHQPNcV8qALbFKIr8mIYvnxKz3Y6AvXlj5IfY
eSuCV7SCNztLfQ/8Fw8pE6lqWSbhJV4P/xiGTx+crrSMr+lqEh6xs5AFm0NvAyBiaIuw/fG6bvwP
Z7D5UtNBuR44Q5TmrsWWpf4g9pbFQpeNEoFoHvpwtsCb5HZ2RGzbO+Bq82j57rSmNneQC/Sbe4Cc
tZv0XrG4orBkS2o9tel/smDyIqKfXyYY3f0Ql0HtK1i8ubLHeYCWm79X8mzigWYa8ll98m5QNFU5
KG66lV+N2d9UyKCTpzCKfTamJ2XuQR5SoXuHiC3eygQgdtt2VfuhRGpqLDR4j5+iv22oV5b95kIH
FqrZjoCG72tBKkjWks0LU3UVNaFyAgcKfXiILS3R3/kdFKiDi2E2LXtCL961ncLE2Qt+4R+StOX3
WEXoBtD+vWQUfjRQ9qBT2VWx5DiA6lBiSphdbz7efUv36AOpuv81a5+FJSLWxBvzNiUg0/RF/Fgc
hnQw9y3poOJ2Xdmaot1FzWC02QqQZmo8PFEBUIjJjf2kEeec4h5OMX5mieYXXalQB6/FrvVUTfNw
nqZ4fkG8vl/c5uSpie+N+T8mFCCRisVbWS5t4oZDDjqM5CiiER8FaNANIzBYTHh3S/FTnQsMifvA
ACnkPp4UUFYjhg0azuFLufaOAgbDyEWfbVyCiVvaV32xx/o7kMgK19j0PNEkyhBoh53rxA/vOlNp
TYJtLc4AmzLbwQnAyTEoTrQFG5F8pxqFXKJjBstDTYTL7iO+CMjo3tE5mbgcBvNNPsUrcrS/v82C
FjEHgwFohVX+pa3CiPq1SEPEUasRigN8heRRQWeX4Rh6mThTHJvWt8Prq+ehoJJ8ujwGWBVftcX4
FLUjRyAk2VGw/2MQgHB2bfp2skKzMbK4UQK0SpHA7VhA5CYiaMoyHpLaJpcaABBI9pCodfEVG1Yx
IbfjzPZkSQU04+gKg7dXbB1ExvxVw/sl1m0NkMS/pNJvAfyqr2gr3DopAtA1DNPb66Hla0KT6pWB
j80/dm2PDpt9ML7+HPNy3UrSDp4jDRm/m9p0W6PUrLG8CorHW3EshUJ0s2DTxviRhCzO0aXoGFX6
bczMFij0Gox7t7x4404rE5Us+t3MToEXuv7NFd8w465rptObuWDcCxQOiXrVOaTY5ZZpt5rE8Af+
+ETgIkPi2LQE2Ioo4UcH/4HIJY9wp3JBmRpQTniXb2DNeZswvVhQxvkF7eIZXuoAh6l/GrC+u6i4
CWZqtwJVruEIiwNiFGKEJhJ1jUxNLKWodDtkTxTSXYDYFW1FRUmp9kT9vnijVtRwdXkK0X3NhEG0
3YDDRJHMmN6u8SmZlphcReL0H2E0nO4Mlc6cSleLB6lXyF9sbKSORiamGRnwGCfecgFwdWbPep8J
yF2owbmtjVI7o+1/uR8up6SvTowtwStixDGa6QT2oNAq9UOtw2DrAqvRnGxP2PFO/uXjUi8RX1PQ
50lb/xN+iRa9Q4AKVIPIzHuN5YjyZFlu178kJh/OUljeFHKtCk/uddH0iSESjVyi1VGgT7f0qucc
3cQh1e+zjcGGPNGrIyK+f2WqeXef+dS3CzelwLJPUlFu3BSHt5aoEprlkvJIGVv6FgjcWminCjBH
RZRU+kHHs89xb0/x5C4g6F/a8hwEb6kEA/rOO0QA3U2pE5dytnLxYDy91yX5MSM9qGmr2vnsSmay
ol4LA24i7L+IQW2eRhcFMp3m00eHVFzQG5288/6NnAM/zgtdHcwUIUTpQt7GnqH6Kq5ypRbHTdiD
g7/g/lv8YPiDkk0Ow54kqdAueCfnlydrJr7uFbmF1qFVWcfjZt8nlCip+wAwoEkvlSQJEW8kx8iu
kSmTolaBMVoK8iVI5m0RQlL4YOCyiDcmbNRw/ET08g1GFH/ARwGRqGhDF9/3PbOhc6n6ksiP6m+w
vShkLm0Fhx0Yvw88slZ0uUPe7nUsvdC70KlaZXmKnjkx2Rrs3px3cxHxNbdlhqxxJ+up0vMR1tC6
M9Oya3Hwsqw1GrDpDmMT9Ejoeas7+IFJ6/5IVQ+A6U2CbyO9gtqa+/K7taMir7v0SpXkk0GYCSLg
8eLkqqMMKibWeUsIRUhCr5010muqCdXE8QtDLjrvsXiDADuW3xT22WEGtLutCjhGrY3E/33Byj6y
oJXknl92zdfHg4aBFxDWZMeWh+5bRxdH+Xo+w5WsCDPy9mofBiHs0DDjkPKYUjC97kN02IhEmIAr
oTNpqoTGndCE3y3SVgN7caMGGVNXInOaKraLoWkhX1UGjHDtX1YIdJBQyt6XzitdJlS4EeZ+iuvQ
mL18jBJqq879cMpEM/VZksj9ggiGE+nvSoNdB+hm72Vn652SLDpPRmq5pjpm9Jh5hXpVwC66zSxb
XMjPtxRXKqQWJynWx9BaOR6Tv/qqox50pS8N93iqDM2gVQyVxi8hAKakJ4iJKfSx6eu+go3A1txf
x2BTlDU6Q892LvkV1v2GXiVakwQkPL4T/ZMC0cn6v432BDXK9ZvlYaM1H3YS5zgY7XQYdncFYQld
tHDrg4hdTzWnKE9PDI7Qx700D5LIkRj2B+uRLeTWet4o+Dm88kBVp4ETwVdt9sqUS6oP4Y+7TTZ5
v5gtuy3m/qEDybMMKulDGKQmdwdRPK8uHf1q/zc4S7h/by0kam/CxRD1zCLybA4fUQZ8Lw8Psx+q
ugtq5XZ6KTUDNI05xtG23ja3avUwUEqzxlO7gCpWU7U5pwphR0a3UzF1mDU9EUXdxhHJPGvUgaqr
NtpignUCkJs95lWJliK3DB2YcpC18xStZ3OfWqHiiCCw6lxS5SUl23MsLP85n0Jj74r682CPnCix
/2X/U44ijaASgXyvROEaH7Rn4ETDFhIz9rh5nT2UIY24tHiC2glHHWtGrft4Pz3rET+b5qG3D20W
5EAhMurOF2syo0amzvEtLF3LZF3rH9GJZk6h8skAvkkBpEA/FFLwqGX7mWFMjSXGZznFJiDOi+ft
UoZqzZoQgrdJ5ZJl27tKpzlC121ByriVBpa75FmKIPl9xN8etMC/ddA+72lp2YRQ1ryne/eT8bIr
4Daa7GJHNCoFhh1k4cnu+iZEG+Y5Op/2DxLOmizeXyfjme285GDPrJYpib8c0A0QiMuNB+kFO67R
pP2W10dpc/15zFTmy2iV5WYNLb91TVOhOizGxI/KgeeY7WonS4SLkNHXaTtrdLkkVFPursrMuQu5
9HptHPXnDLQ/t0pPXNitTZ0lgwkLGpvyHICvDkrTO1LmyOHQpM7ubg/g8EdIgZGzAzUJYbge2w4K
VFW1NA1E4AE8a/oWHOOtEbCwOSU1VcwK1eI4aN8xunWA0pedxs99g5khFj9eGi9+XLDGj4RKsa0T
bf09GsPLhkGKrRhhyYLLBFmS1HEUuoTyXCKx9yCWTjRZ9qwDEm5GJDlrCMVCxQEsO/WDE/M5b2w2
XIDGEwPL/VVd+t/J5uPtaK7+n/g4Bs+zGkX59dQ6xbAazXidDPCgZBlFLufiM2+kysj2TveNxuWl
ke/qCRPiD76DO9hfTCTY2GnA45OekkxiGGcZIFI9DrQQZYhNRAk801+679pfiUoE8e1fVxHPFmg7
u8J4vLlDNmlKAp6+kSin9BEZDr3RGjXvIx3iemWXZsk7L5uCkJLm00k7T3GkJFdbWjdhmPzsm3VO
RMMRR23p49+H57DPnr4DOGt561+oKPEiJTcoFzQk9qdpwh1fWpGoMfYyJx1Rqj1mj2wBb6FZIpLL
aMTiKrArk0bOd9QMJXxRpjzw9/ka7Wf0RwH1AXfoBczsi1otFdfTVyX7QkVIv69VabfH9F2PXcBu
94D9a/swqtrwqpSqzKBCKmcB/7v24DkH1exnsSBJua+3LZ4NxyhFeCLirRXS6kUH7KFTqbCbBF+q
xJUBrXAEUprg8kOSczRGh2OrGK0bffJjevC+CSdlI04FVGezeeeNbKiGtVzFFolpwLpk7pR7hFWG
ShYP7i/IZWuFkssv7Tq9ALpeRG/BtWpDGmsGYPi/mn5BuWmfoseSPMCO49staKOzvPwXAGUxj4Hy
KnsK+4j8H7aDAn+OcNvjJsJUJqf62UHRowCauELBQqW2XASXGSRUOHQHSiuSOIdOlYBOIQFcNEKa
WDl6GCrBw5EWvghEXmo1z8C2n4t4gGeTLsDHshjuCPD7L2M1BtEotDm/Gd+cHuYsKR5YbzXYahkU
6Mwx68yRbU1lAjdBe2q9muUsv9Ra55L2gTQZIApJZYoYn4GkVvUOcf29Gm5TS1ApEQd6dqMipogL
0Bceca4tWBT4VgpRTwDmz2NDbomTpx4wUut7pdYw+DBDCWl34lAEVQxdFX8e0mq4BTIRMPs1SH5M
qkgOAtP/CJ1qNbpW2qAJC8dP95zMb7+sloH+vppmJVt/NAuqGr3yKDs5fK8Ls0PMDk3J9XU8Y9JR
jJvlfKb+YnYH8pb57m3QcX3pN7mh0qp5qSPPfz5Lv+RYzQd0b66n/vd/nbSg8t77jkbnMAICWLYv
j0nHIQLnWl16130vpCQ4r8lgw7NE79uvkKHQGTSm+smzVeSfKEXWd3jlbxubfQUctnYfnF5Dmrgy
vSxH22qf4JYkeMPVROaWBo4+cdVNnfHVrfyxS3dmNc3p/Ocgjctc+vUdjlgvau3/xZTSxLeQIpWK
gePfSSjNCwsb0p1aT2HDnfUBjtBV7vO/qee70Nk3KMUWZfcmKV8hkeGE2UNWLi2CxHinxJ6cWtyf
B4URCjKGavXLoSZf6b+ucOCz9D8zk2qTZEkXGB4RmtIZKtEBYMu8zKNYyPvwaMNwGQBrss2hodjT
+zznbtbK+ymPQ19qz18BKm2wfBrJJltZyk6XBj9xixkkEo3OyDLM/6LflbhVX/KcMaRPljlpMgV+
N2uEU1fl0OBZP3YCUTBhtGYJ3Zo4PL4huWAMcgNfI3XtDgGY+6lQP5bJ1wMB7aD4AvkNtMz4g6jk
IZrl4DAmoK34LtLvkoi6/GxXWE5InM7m+hhEtA7KUil1xR2HDK+WoAtXwmLJ0H7ilvz/2Ra9mVdB
7fqW3wfg49sCbZ74+E1N2cigLupWMhB26AXjcw5JRoIKksvbDqfxhEiHtINSLqsO32YvnvGWEzVv
WUOWnNsbNJnn0/ezlm7gkjYmz0zm2vIFo8+9c4RR7Aea4mP/UunXzmSfmptJk4UfqZSR65UuC8Yo
/lCJtmlg8NREqApGawKNlX/k1GH/Xsqsz+ABYBKV1zLgjINMZvknIc41cpEG5SPJuWHfyRSl2/OA
46Ndbp2k9OieHn6gQ5HtlWdgFWVjzDnBNr16yRW5dtFtZHfUZnxrewe7LLm8nXdgCo/mUhE8dqXF
qB8ZuyQRBFR4GOLFFe/inloAgsMiJ8MWO7vl1xmfHyLEKzkIb9fUTLxpo8OlxDAsah/sm6Y0nIM7
V6eL/cc6N++Ufm4os/BSJle+uJ+pu2P1t6ngtRVeAeeEOcFoSLz9GwIueqnjUiqgLIWu5wYggLbb
rI5qWH7H3fIqllp+J0cfSvawPraYV0//+c+sj8f4Bjk91VMUDgaCgnP/SbDSeVqUouHpdYNtEeZD
O6m8LG3KnRNXOfPsN1hn1nvuwd69zADvsP2uq1bDf1MwAxbXSUExyfctKqBsLQfjMWuJ5SVnkwoL
NGcawtooQ/TJDYJD63DRQnHlg8IxeB1g5VIBOKwoHXC8sKL+vWY1dPC4l5KBzp/Xe9onS1IrEQgM
QJajEURavLhnzbe6FvnY1cRW6i3XlB4KbydAiJQEaqtaSZQ/OM/XeyndaD4/6J/u4KGTh1Vc5Iyk
VnbPz/NwDGOa//KcQknET9hqy9+xa7GLE/zKZtWtLLZ7yqPfpsx/vg1ArvI45WWeq6+oRs2OGrft
8J+NRGHQXQZnDzWr3xyN7hUqkDqGq5v/6Cwd6sI5oAUce3uqy1zct0z2h6oNMapiVv8mIsTonl23
jvkTia06/84AeQEcW4voH8ny487xoKKkqYoSpSVkXaNO/SG+MurdVjsvliGIckcEM0iFXgFGXLBK
2h1ZO7Uu+6vkpoJDSMBnznRY/rcOSM0un1NWBY39Tt+XWWCzE9qlmINP7ty9UR7FjMyC18xN4vuK
A0X5PZ1pHEK2756ZUffCAKkt/M8iYoTW4dmrzAdcUMMTpdbGk1mb4NqF+DcVWK3M6TiDylJhhG+6
qhik9EIzGSDFwBFeJZZZo+SQfLl144Nebm64UAcBytSE5yNCsymSZcS8aGbQUTcgwYzT+6pbD167
kAeMOOHfwM3LUB88IRtPilksvSHv2zTgvWaVfrvuhOywFO1BPoeqoq8SFyrDzVEzRgTIJ9Wn430K
aRkB/o1yBg9UnQFw7TVaUjoZxSZkkjhdnJj7+UgOFT2G8fOx60QCUEF0cK71S2RzB9gDgn2YSPjH
0orvuuM2BEMiVNTMvcjtVjn6jgk4TDmH3U8eYwruRX9sfcJZzuroWeW+VjhkQi5qDV7wZWKmhRJ2
OddMBrhGn3QLDPXXVbOYbJlbG94r5DVJG3bDqNMkJBD3NcJnM791kRh2a5x8XvEc8LwQuCpQprmz
zLdhcj+S1hiX+CnODcTDJohK0vLkGH1ml+1+VCxv3HaovMytA50n1BqreIJsBjgQApp2abYjco6z
Qa8UC21+tnE7kXnqFELlm4AWnfHNNNlSx5h9bGP3lyivEH7SHwbPUiJOHtAu02MMyOGDe9RJ+MPg
u7XNKIZfuhO9GxqMk2AzU8iQzCKJSHYtn/XwqIQKeCeyfEfy7Wz5jskOC1S1Tgj772MngpHtXl0h
1k1vjIT1p7aN2JQvl+rC4VndppUDZ0TkrEODuRxn8bOMq0Yftmgx9FkumlB4yR2sBinRbuBirYFV
iADi8az4gZYwxES17qnHqbZvebXBep10eM3Hf+FB/whWg2PFi28Gq1W69EeFDsaMGdW3Ri3Ak2HZ
WFKhnlyK1qDKIxmnPQo7YscUaoSGr6iBRGa3o0yHM3C4xO91Zrq9tEgICr3oDRUYHDiyArQjqZCU
ccgAeZfIx8LSRJZXGdEx5iaA2gr0/MeuJAmVydA8/Fca/1WxA5gLhVR0TFRICcFl40a83bSx9F7C
2ipWAHleOJHtU1JdaxAGJcXWfQ58W+elY3dNeN9YQ30mC6eo4g4sNTJh6sJx+fCPpzcvZoopJeN8
2DzEGziwlQrdqZBE2pO4CoBKbAg/udmSVOvOTw74YAWDIFyTPZrVxLa5DHROxU4FHcn1L3+q+bt/
jvprJWyFCEO9CTuwycXrHKYOEZaXmiZFp3NVRpb32Gvl+2RpTy3NKxVr51ffx2JFPEYXCx95oaoQ
e+rQv2Uqr1fVFw3rlmiG2x9gkt5u5+PoOCbuK1gKiqUlK0EmjLMxA0lMWYfACU726SZTmcZNRTuD
3o4cRWPILmGexWVTAHQVscPm/FGG38hLIWeITJl8rsO2+lRPl2CYBbOCbOO1fQsncCMiWdvhqONW
P10lA1yUZZ/2ozJsSNz1x4TA6nao8RhVU/GX6i4ZZCa4uMafwHFIG37aNgJvrwUPSUX95yhRSfNL
Rw6kFIr8/ALYWkSuuvwScH7iWoioKayoWWzRdgQUwNZsMbBO0qNhwuSf3q6AP5VQzjqQZQYObEN1
Zjfgj2lw5do8ZD6ZHiBKn3ydlkn0koQQLVTnInJUY/jkPM6+QhpZWBqY/pN61McPd+kjyNR66qPg
D0pLwYOs3c2tsS9rYTZp/pM0EMVA81bmMtZrd48azwrInk8aqNNPuZ5gCdVK/YwV+JUX6LK3ffSs
njAFzB9Wu/Fw+3QupAbP/prOo4RX/Rm3Ctunr9+oc05slkF9875F23ZGIxTyjwWYzKePRf11eker
Xp7v72jZbGxEKMD/XrEBoo4T5zdL3xYmp6JQmKfDmDuXcD0hmtU4PV8Nge69ACzyXiD4m/4BdrBJ
m6WspaGln5v1vNOmB7HUnd3uP3G4GM25j8HfQNuWpGMWbJ/seP5MkbQuxigB4vRXN9hH2tbv7tjp
laDpuZJCYpFtAB6TfjAWxBNo1+SR2HaKRpjyY67plk3JA5Xu+C+qg2zC42mwhR6DNriZt5gAwnwr
27Hj7dyoa/dF4+yh+5UB87b1GEeMhBBoVsAeT8w8piTNteRqlSZAi9oQE1/vxtYgPzxPuNXVy50S
VSLm4X2jZQWCDl1TqXkWuB9zB5gq47WWdKNKIx82FaOWsVcJxiRqGAkDZk/OqyN7jUCkeU6j8NAj
rBdnA2XmIRqNpO7Iqz2PZ2OYeAm9b4dfYHKeKsqPB6Qq5qjqbTw+FFdfMGsqY3tpkzHo/E0yphic
PTfIpmyjPd69Pewtvi/UESgTxIzNzBrIdxOqGTtSnDGCAI97l39+dsVZpsK7c8sgkA63kduwaBsU
+mIW3wxiEQztmjd601EnT7Z45CRe6DtnitAlZg+Y0++FLJbe2NhsqEn0vJT1sFwvCjj5XqefdrMW
XQFKNW17ksYFPq4vTZZj+X1EsNEPYrBL8EFb9b9n7zziVl1ev5dWGp9ICnzmKG0mZDoswuQBlZ5S
XzN/T14JOhgeKKp3dRtzg4h/oRjXNZzUftVAJFqKjC2eowjpubEh97uzdIYQD1+dEelsD+X+duD1
vomixPioWjqYQUhJCGqJT/tdns1ofF9Uqr2Xwac4c3cT0yY2w4Ng+eR+UbBTRKy5RFypWqvn24rm
WhSnFaLfo3EYYcmowpcNeH4gMIrzkfwNmUCjkNl6AbAZ+6OonK3En72vkMApy8Pm1GcHHtPc/BLG
z9tTn/WZNJVe1TK1EjXi/PxNgg4EMCYSiaANY2UCdoGY0ZLdwNxMBpjPWvhkDSBAolOYPDN4Xm2D
rSi2FgS/kppKJ4Fklgnt8ZZ/2hhrvj0WbIvCAKP/XlBtVks/dL2IpyEvAcZoyJYk5e9UA+OEWoOA
dAN4TOnFXupvVeqzeSHRxZUEl1YwA8ajH40oAfUr5UWvW23iuUzvlTDlRj5GjlqrRe/PYs0mzgis
quKWldxaFlVPnYcSs3yPXRIbA35SDeIXCBpvHkIjsdYoXt2KL6sqFjnmpX1K2eaMokxcaOb47wV6
TXCQSz7plKPVkHC956Hil9nuQb95m5EI5m7Cp4WFLgT8eH/gIu8ivhl6qnyWvjp+BPjXqsO/keFI
g8EipX1MGjvBIQXXgAgoZEybskO3ye3/M9TW+ybKVBkGJ8wr1lde6C8xkUL2tFmjaSIh0e1PXT+6
8Cnt9fPLScllEV4xhHSZy0g43nemDv97Zw6PB8yWqg++XKSo8u9rHNIy1KVAIkxL9D2PpwVZceSF
uOx9Wj75Ya8acW/wndYyJH6Gy/+OtQsXgmPI3wZ688QlOAH4GB0sjcOQwMjesHZIpW2KAnj0EY81
AxsI95y52c0xk/QpLZHpdcuoNZGiiW/WLg8TR4DZX6xbjglxwRcma6HUOuotvOMsHTjTPEPv7rRO
HyUd/8TjldFAab6B8jylyRi9ifevf/8NNuExOtD0gSMiniVjNAJAH/UzzAPIGEXPE3K78aJgMHQn
G7GenQvoUZ9MwKbe7g+rNlHsaWzk9q0GlpY6HcfKThDClX2VnwxSPmhRXSgtT602BwG8Wat7N5bj
QyP5HI35R4OhkvdmV9NPLXf+0tMosEn+b3gqQZoY1X5XhDOx0M0fAfWVHhzTjEgVB5ZLY0ewbPgG
otMDqeckuneCQWRzMFqbLbf8MIAyZ9FBjit/+h4XTFSapmgbPPrBX0a5MPZSqAvgjXz+/krIH1Yo
cizzlscekvhpIE2+HXlJpwZRuoBmaTCeHsDJq3vLtCr1uygqPlVYqnDp5SUMcCfnU2B458iKPwH/
Obb9O17KjNziGlUcvyZN1M5/nW1wynPv5vwtP7BEsI05wBl0Wj/yCtIaNhbRT69n3iSEHfBDQ3YD
jBqqwwg2yH4e8RqWoog8OClS0gDj/ZaCur21r0f29mQtIOafNQNWle1RnGIK2Bzf+mUTrr/rPD8W
RAffEtCiIeTjz5dXkKYkJhsAHb4O5VrDoPVCcAwUKJGwesALyFqKETEU57JY0Jgz+AmK6YEzhsbF
k/D69Jkq+5YJsFGHDVrS2xsCzduEPG6OpR4X/18G3NjmIMr1ouMZMX3dQ0gEMXQMpw2O22EIyfvv
4a81kwv4//BDYQaCYUAuAt+cqtJGwfvodOPLKB4jwlH1t5EEXm3GyZ2PtHIGPbxzmVkPYP69OdWV
QT2HXPdt/zUYw9Kvi6PvQ5xFHEgILkWq1B2YR3cQaUZBDaloyqDeECHN0VLkGwPEVjijN/wOfz/A
e60jPpz8myeZ+hMdsXI07CYcFuiLfQKgK/YzPgvff0kWtL19vilONwruxEZpst4LfBtg2traZY1Q
7lgOiPyzOlpf9iTk35EIftGGQH3Wg6yA2oLf1LtI3zBSfphdB9gKlq4EG/RpuP0MhYi6a7aJ/WY6
f0INHXqaIBrbByCYirlyDW4Oq65cjVK84MElOZzaWZIAExBM3Bl7ORCXlXy9nlkzG8gdL32n4K+C
orRKlYPSh11+7X/kM2dgJvyS/WkhgeeAUlgkR+AY4Ru3lf4SOaeMd3gKGG0JeC2i3MOz3+6iKVJK
gRnZQJ7+4jCJzJt2SJNEX8SoEn4KByP0EcEXowT1XpsxyN+5R2Z0lkfi1SwZOYqbAPL0EReBCLSb
CWtlQPjRRrQakUREkwQ3NIjI2osV20Nl7J8yX/KxL8pQ7sH6+HsCHPmIrXGhnW6Yoh3XZxxiApBR
FbFUJG5r5MwsrfUFAFYedB6L6BlIycCnB0m0U57uT6/ZsfgoV96uMqBCzj+AT0x3GtrJHuned8A7
aZKnSTDZbJOc0/mHQlqTqUQgqxmXzJlWOPSJ9R1Hu6zEvYyMWDsxl0OxpQrZ8ee+HGoeBNpEUei7
CtvsLSK9pK0tGK/5SMPFta1C9ue8PZkWvDPCSUtWLmBCas6J6vLyo+jIyMWXkLZIkiVjlR/nz4ge
UhsnbDaVKuHy7eMm2UbM88IjCxQy8NkdJAwHFPlGQjjPxTs078MSzbBKch9Kr2H+q3Ghv7OSGWSM
uDXJc2qGP9Jv2JWbovXkAWGFwh2GDiIRGMlNZkCCcJNXV0OeDYQ203D7J4CRmQxk2p7cJIzMXOW8
ziFP7Iv1GQG/dyS4j8Xmx/w3QMlqlvDZtazR41Ol2qbfSSZRjiYyBiQXYWdzj5JFF1BM9b90EVmU
XTO+R0cqIY8xrR/tqUZnh7cMbKsK4Xylg4iIktI1KEsa+CqcG0Lmwppin7LoSobHCsjLz9opK7Hu
Kih9dN4cGGV5ZO+xsRvslSoFi2vC/EFaQx5ugYKFSYdA6QbmTlWUAKh1zjZ6czQ3UPUx9s4AsQZE
N95jNJgZ1ER9JiRjPOP5npW5W52osZFo2Wt2i0gSY9SiPnzvAb1Q94GwwYuzk6PalO9JGMlz+McX
4I6xIWMagRHD8YEsh42UpbcBIFw7mOfG3an1LiWKTnAXQy8uokaQKmIVAClLXKW57tP077OnTy6G
ObLoG501gH+M15Y6EmgwlQ4bGLQ2K8iRJmLLEK8PUx9Ny64bx5aE/+5kc5KJkqG2/8HPjHY0Cs7x
YK46GbvblknYjOFTSEru9Eq47SwE05YQ6ZF4/GkZAtoFuC3tKlXQ8DmD/Bhk2SXc/waSfrZk0aa7
QYK+0bov3OR71FWxZFJBP/luuUuAn6zPZZYCQTe79pYj+H/c8svVwG5FQAE0juXY+/MMOWCyUr/g
MuqHVFBq8VNcvF1w9Eu7VR2Pm5ukAoaM672U8XouGbt8QUBtKj/BH09M6ADmh5iyq06/9a3WmWd7
4JhG8sml/ZA5auhiqzG8tE7b7lq0f6zqTRh5YU73wlBShy0xYoXBPX6sIfWnL93FTGQWIsMf2FuF
n9VRuCnRzD8rm1lhdfGNIQ6NjobpVlS0kBJowCrKNhLVOO+h+S5REOL0uGPVWMMmJZod5RE7Zsg+
fPgk+T19aQdpT2TC3wODFHByuaNmkIjvpvApybCnZQ+leoSc0Bz9P3yiWFazHXAJ7nXIESBn1eo3
KsuidFuw40ySGhIc3qg1RvR/EaSeMg75w969AtuBa7sZ3eckoU9k4/8Ch4QeFfoHGPZ+FSYVFIY9
CcysEmctNd8MMGELY5il1fryM3LT3UZ4m0cWvnX3IY8oda7kAHU0PQJrKmMR0+kqzOGNopKhVQA9
HKD73S8FYaDiBJY4mZBEWvCkthbn9pBWy9AR+qOVO/tHVnsXzLzuINb1EHRLUasemaW+Q9fDN4Mo
FiouC7HSaQ/6gXNzYiZRe5VI27Ino/Jmqfa16rSZHgXRxHiyvuy3QsQ7iOwuKyPx2hw0DVgOIuRj
TndlqW7gIKFfjlRNDqMy0oBuNwb6JCGvaPPWNJtz6tUJDSqNnFAgOoBNXL1rCqeRei0oTNzw/UKP
rpToKmsiZoUu/RMz7LMVbh0K4qRzloSMXVQItUfKAEhaQH6hz9SgYBJJpZC8UCyz/NWx8+qRB3DV
s6/C1BZ9zCyQE49kQbbCubGT5iso1tC5SDqVR97PumUC1RrUzHu0gHg2rvYAU5B3T8UrkkdWCFHQ
hb+CCWPIt6eOd85xjvpzaDdo/tw6rlRcfoVwuVeRr564YVwuSD61ly5DYN9KiE26t/C8n/vmy2oH
qpEAKz4W5D9sK9CPkplyNlQVJNOyg/ozoqA4+f5f00PTRgJpLP3tqA8/Nh760rQKpyiETQKcOJ0h
YlGBMaMmx8BXapV8sD7Y3W1cU/SnOxHuX7FoYFp6MALY9PNGuJ4J86tmXL69ER/1EJQApNWpX76k
aIF3Q86dbfoEwx7X0XjGzeRdGGMXuKW2uJG0c8Df5n+G3wGG6SlUnXQS7sCocv3n38PQLUBgqH+F
ucZLYd3rgc5gZuFAHn+6FDXgGv3ODjOFU7xI4GH0U9LMLjWfzGc3Pq4b/EiX9+hCZVMR9/EUDyAA
IxIbHfePMvg5U2gYYGUdWEP1e9Lk7Lm5ucgtguJhvhiOyRZxsIxYVVJXmM8XKlV/LT/9gETTyIGk
w/QCvZ9wqXQ0FJCiKTvLOHjpFFAoZZaAj1dJPKEyK4A3SncT6VnNuJroT8Woz4MxHo4q7UW8AmGu
ASPDEg8f6+orQwm/5r4P6gcr6UDyYCVoFd2VPjdvi02OsMawiepmZqZGU2UtuwxC7c+YjBDwGZVT
7ocffR5EJpPZq9XY+29rRPL2dRnrTo2XkB0+a7KlU0RE7rAyvijaoIIWA1Ynv9V0aIzT9AM2qYze
0jkD7ijqCtVoeecIn2EQy+bEqDZmx/PkpzT0+RWZuyTv4sCmGLVFYt1yHAzqqUZC7ElF6B5Du38G
P3ZUEApVLBNOZ9vBYD53arWFj74JvtP9EoRX7/+2iHdTBba6IA9EdewmCCcleGNd3DbYPWX0Gt2s
3zyyIE84FuIM+HNwuodSYmy85m3LM5soEccNr+ExiQGMjv/yZtxHJ/37m/ycZfc76Zw3f8ufZJvN
lmK+NbcS+J4Jf8XgdwgZf4hsrz8+U80CHIUCXscUYf+WJc55ol6FXK1nnFl6k3+CQNA6RsXbfwc2
6BO87KAP/tcrlv0D+m06YeswYbw9uOJR4NKirNVknRryjMfH7TGX9N8zWR7MQoy96f5Be6JLSWqT
1WgjkIXpXZGNWA52nO6PvNbFUBu9cr2V94NQZTA5BSBU2wrJZ+MQKxDhCRGxFW82nmzDrPj90CS9
bdTpB7suEQrYizwSNMXO1INNxZtbQ82Dg03bCmiLPrfdVhR4tJktwZZ5V1mtHlbwjZSTEPP124BK
cQWDEa3a54N6roXZ17XIzA9y3Qkea3/Yt/M9cNuHwZeHGfuVR1O12tjYse9C0fX7aZoKPaXe7gZV
CtmDC0Kn/qiL9cv3UPAtB3PXyN4aDs0dvAKyKIo4d78byP6A58Od29NQhDdEJCyxjxD3rTkMyQvj
/Gx/iejMsKZpiUIboIu81lvHpcP9iTMhIdIlvBC4BCgV9+P0yUTxI4Ys2lSJZlxRoNiW08ZqDwGQ
iJFb+KtXTaozzgXoeK23Y0O2CQnuYBS/tsei+QB7uc2MnQqZzpwvnEu6rPNxDmFXxGw7eFKAHaGU
jws0S2zWZblEgU2sU9hFZ79BOzFY0c+P739fIvofAzwXnpPOPD2oU4ddI5RtEXmcEVIQSBT+kTuI
xv0eskqaqrHepR7n3zL7XUMRfD1o7HmknmOUAUB1EjqgfeG5u8HFA6xa1+6Pw+5uCx2PChKrcYk7
cevrTfr8MjmW0z9h4XDAz7znh2KFQ50OwQVth0jVux0ml45i03Q2sJb70pBcCZraCsoB0YNUI1QU
PfRYJzHaqs/vTtXwnTPECsomWl8jIWoUgqFcMd0PpifQD4764aeAzliW8NoYUpCKq+al4+UlPmK2
x9nG553tP3T20Ehk4/KeR6Fg7UqmNneL4Osw88onD1ga1EYl8N1r8sP1jvcnZQ8BtBpR7leDJwMX
kq7V1EuQ/fq75ptx/aYhSPdefeLqizIITvJVmnzSFtTpvWTUxDO0Gwt65v3vgCIs5C8Rxed0epEL
sbp+8/edpRp4XTwJVAXKhQZRQ0kqQr8sSOdn0DtkuQLsB8SMxGj9FS1lHWt1BnbC9UnzkP9edlCi
0vq4R1ePxusv5QtWbuc4F8kmJh7AysgeKGkBsNDKak2nmOOP/eZuL03kOuB7l/ZFFuJSzIKqso0F
q2YpfzL5NNYDt3xfLi+aogsNDjWZUzgb8ELOwO+oDqV5mZunQn75p0CdqczzSa4nNlk912K+2Mde
TPbMd+6I2drogq36bnqnydqe2nK8fzGzHPElCsCkzXXIvEmjvrC5S4VEcdMjX0HArss+F4SzysKt
0UUfVz+T1oHFGExEpQa+vKV8SnwlRKh10KgCt2k1z2mj0wJ8LQxV+qMZjJTKgL4fWQ7teEFXXyrn
VwtjSDrQh3P4tuh/70XvZCFU7pKpDd+/Z/ckiJjqRdATDlTx6PFfIRNowgfbUZqoq1JqPlUk8uli
660AGU8+AS01zKi1wOHvoSJLya8SRfr9le0HhhALurGGDNpRIfFNJs7EI1s5xQLFCEJashdpXdZb
Y0VSzF4Z4Dt0pNtfacyofmFDk5C2nqVgX0IrtsLhPmXGxUyl/yWQc6AVC/PKO+tjkFBNHAZ16jRk
aZveYIqi+7lTKGDfZzoRDo2WG9oWcqM7egAA1GZ4n2Fz6ZXcZAZ1NQ2TNWsJWEyJ00Z8GiJ07ajV
/MiIoVBAqs+ZvLKapVTjFinJmRvlQeyTc3ve6mLkPHCHThcvo/r77preslbAO4wLbKktWrwglRzZ
M7wgGHhJcUhcCo434TwpPS+N2hYtCmZJhvmC1BFluY88u2xy0Idnzozr8DfVjciYzBwUuWCHDvYI
LoGk6NrOQjC5MoaxOUmKo873QoBGuEM3KK7Z0xfpjFyQA6ttOk3E9wkKz/dj5XM+cGZsxJ4MDiFb
21UANke7pxh6D/5pVNn4D196JHGkLlyAdQitP0+YBZKZVgv5qA2RVu+GrLdOglASHKE31KkeJoJA
Wp8bg0syuAnb7fKcj95DnSQF1yDsvDcve63XYLo2plYQi/+tWY8ZxUBvMtcjZYI5f92p3yMYpXPt
ByT3je5M1R1cW8+QN/gDPmZHIWHOlXsh1RpgITkjwgOvdHlJo4l6JzT+yrX3RCpfzSfbAmKyZjtG
IvT3jijzUtsQJdHEduE9ltxDTbNQ0c3Ut0OezyLmXmwF4WVEu0gJTpXokpi7LV3JNO6pw78B3gIu
/Tq1m4XjoEcMVPPt/FE7apoE45YWJpLA3BNFrew9MLA96RJoHIYA15Q/fFe5gK5n12hobkQQd+tI
/D3y8rmwzd0VMev8Qi+nIw04ibwAbxIQrPPAm+pIk0W2iyU3kE50Fo3CLZZftzkNUGD+ugRq5HL8
xmwcNU5CHBgzFRaHnqy+qlUyL6tuyjTS7cWci99wNaFwBHxqTeqzrwFPZyfl7LKUjAHsYnRZiXLB
iYhDM+KWwSu0YbcXD8ew7yawvV8ZYxKxvxE18b1msDAlDWF2O6joOEUzBYhBvKXvkTUNnavNmdTp
xM7c6jRTVXOOJCZPvujl+xBVr3x3czWg1X3+iTyvxpLW1e8uUG/Y4oPHIgjAz6RBrzdXwA0a9HJ6
MIGsfNeSf8lYVNWAomYF+aOr8nGzjfUvYJErcs5AANRk8yJyoNn+qfJn4AOPGgfg2Jw8xOnvDbIo
gR/xfW1VK3RU787SAJZkvbzxZARqwWXz2xN8qkhiX96gcvX701SfzJLWs9d8x+UFHU9iaCotwf0I
Enw5XCe9b2mA7nbrG6yZ12mr0ceUgO2zGyywROs6tclHS2ef/Io3b9Rn6a7kdOLi+iYh7dnwrerg
Lu5COBmvR1lj6ihYzeLb0TOw7kzFPyU3bAuzA2asEc3pnA2RDweSbgpV+mqNhYs28FlVKfpFoPY7
/KllIKNV6XIJCYDwsoSkKBpdeNgyRkx2bxO4OJX4VEoDjnJ9ST/LkFpy2JEfFEWrfjIlrhul0uIY
wJVK6HtGGRY7TQcgkUNLN1iyUoddyRhf5mU4MVtccH22+ZvO/+6kEetWAoixIPjrF0f9Lc8bxj0O
rGCDp3Vh7IBosesXZ4+BlbaW7qzl14s9R4lOJcELTYDqV46fQ906JY+HZ/ZfeiWVf3ndvdTJpGbb
6KOYaWcBjn2dFF7Y7yR6Kip9vCIZ4fkDgulLtOZKHm6kGHwDG2MA069WDuoY/jN9jPiEOyqIXlYI
NICXb8tgPuxV1oKdcBPdYw0WbEX3yceH6Pg2aznN3AIxRG384fnRzS17KdKZYe3GAIY8wnBN99bs
rszM4GW2hJakl82hGzDvDYye9INwPkXlKJlv6YF1MHPgTHffSqjDsYnVzK5K0rfLAqDX3C/aZO8Q
K+Beg++DW1HUIr8UakB0W1v+GFE147syztYyP/dFJumeJLEn1PdN1XjsbhNVCoeyEKLtjQ6WVCU6
e7wF0k/ADSEc4Aibx0OATrEINziS8TJbVlQSqBLxhtTvG8X4wt+D/kSWR1Mg+XFvbgy3+rKewCmR
t1UKGHvf5As7w5m4KXbfjKstJ6Ui8aAIiAObWdVF2jUHHn9T6aAiMee07/yvxaEyNW+TsnGZ2hw4
NHgi3bGa/kmuX5GccwTeSCLwo/dr9ZNfMDL1O31+RlvBvCTj9UJjD13Zpxro6aDdcrm/g4Z6ACXp
UGM1BV/s2EvoaGPfDA09vfDNre0pCsC8QjzOKbbfOYrkV8DdlGE0l5uJH/KouZH6OYLD7SRH3BGs
uDTpiM3KyE8WrVDTajuoVdChjjWLJ4aEBzcRoX1EEa+QbiCENnjNr5HikVXZHG4FbvKDYr7YwuiD
CiQspcXWS9pyxpXw9C2XkJKeRMbv0PgIAu/O4eYjeAFZga3iV6U6FrNzkyXMcVCqxvbuw2Ha+i3N
w2UPQ9xN/HK1ezTropyvQCGZKEvF8uN1PFpcszvx2hLK5QkNsC+tMaCO84UEKPGNx62nihaNinQE
DjtbmUZWW0rdcq1+V6qDqWo4NPcF4RvIKfVqygtwXoxgXTKA6I6wJHaTUEb3iqBoZEJBqL+VWaBS
inbGXQ2nr+xtJVAes9HEGkXZLH6TYXuyz/yra945FPkRIXLRkyDiaRpBWJ4W8uMP2kv1LLweevA6
YR3bZmyL2A+jPqxmIxkc3bImeqXm6iC0sgDQmD0rtdapJp1CSU7/xn4YP+w2U+MFD7loWzQLROh4
b3MV3EcevVuYy9GVhI64BlVwRBeNni4JZOsOb3b5BgOTjbm0nLBoMw7gImnOFyUN83HZ1/f2eEpy
PpDxFw5hhqWH5aS9aF8lORgp2fxo1Gj36g4bvYVm9igO9i+ci06cugdnpcW6jhdI3swMJF2SjC1+
TFsbjsd+/09u8cN1c1PmhaA3ZhYZQbvIRsGy1xHRthNO5/hnUECRNTEOWuuYgKHm6xRabxqaNary
KKKm5vNJkBJVkKqEbfdvee+WTbyeA0ZuosKGUAX4qE5soAgyAd5UCdQt8A3mNUY69eNLhnbO966h
ehSw3hEYzVimZE5cR0titksrxi7CK1wPxnIoyZ12+cizxl+GzPBD0+4VI0kzaadfvHXw363pHx1B
NCVykJhqJyguEN5Vq2db7sLatBdNOqvVjBVZOEekgVrKviW1uD9xv7Fg/RWJbHkkJ5gDGJRUdmAH
Ytwuin7SWdi0DKOI1xgZutgfKOh9/cjOE5SdVAfE+dWOn58FWlaeJYa23IocsoRnhvoCX4CRpFIv
ZwdCC8QNuyAOVTlHfst5rswKB1y15BQJiflegXN9gO1e98PUOCHTP4S3+ownmWyMBbnSrWTkPEvy
uUotY2LJEvCOK7AIRrtjma1eF9No04DbfHrb2fLxJ5f6NX0onYmNDgvqGqYxyUSGu+g2roHE11Nr
CTHlPG3qkaPp9aSz8SKwN1a0bkQHKrLSL8mVOmXUZAsTD99vEVNlc2TCRGKQVieTbQueFyAcxMK7
35kZDKWLkwEZYm2wWscpjwxV7Msug7ZpY4ofcTPYOnrQZl8wi9v2jY+K/TPRbqCGgDo1q9z0OcTm
O6oP2wrA0O30nXDgkIbWbfevqYphhZwA6P5EkWG5xSAroRENssLt4DrFWEV+t5GsJxWeKG7SDHqq
c2qBLZVdBQCywW9lgg4zVr4ISTSxA303/jN1ftwuAsXJmGNJVKORWdZbNvWtzOTgcAK4nlb3mAg6
rCYeqHAmn/QKOl7LJoU9L/hTbpDZF8eyUPIzgkba2g93Q4ywXi8awhdikGeWu3WrdAuxcs9Uw2ya
Ep8pxtCngFHJtBCWX3F+2SDVZ+hWPNsebL/tZM9t5AXiNKzZbiRJ65/s9mn8zu895hEqMkFEcio0
j+Wt3KSkBeqHlmxQqHanPub+xsPS61VapNK8UJzsV46IoGsJR7OGifu5vhuQl7ycEZIlxBvlEbyf
hgxNdsCXzf0YgBRL2zMeLLK2VAunW++CItuRVc+yr56iseq+/IhsodAanXN2GZplEc0cB4W8v7y7
/pDSEc1qVYiuCSohvWmj4r4kkpl0ETk7TDEgol9d/4wWlnm38moZbAvZKKpDWXKxBZE+ly5qk6R9
zsY66cfoYAUpr6PXDmKAaNwTvw5otsAgwz8Tt+tUDfSKjPxsiosvaw6iUYM93UisKY2DyKDUUR1V
2MV2CO/aTs33aw5OZYrV4hmVGb52dPPduh9YIIP6fGgwiOpseJ3/9v5VkJ8G2KahctBxlMyoj45O
PYeIt2G+mD/h1wmwOxYyDUWcQOo98z13NqmDXA9OGnwLkeYeq6fsHPSQjQmHjAW2BJl07pcwlL+T
vqgW8FDP7oGU0F7Uya/0PlWku0qrAdPN49nYB1kroBXya4TlQnf7jsRQeJy6mvJ9vjHfAXITZsQb
oo8k4ZnoU3wQhpTKKaox80GMatzvGYD89a0AVNYjq9CO3KGDwvSpdQJhJpZQP5yh9gC8ReFNc+e5
Isqyuvu/TQotVnFUK6twXx6wVjyHHx20wUtbV/S2OdSqvQp7fND/Gebe9ZLsNT2FvnO1tnVFaoxG
Ix+rU+hrH5nsXfUHLPYXIECcIo3Ynq3rgVOHS1d/MZ3BruzmAqv+ahQ77d7iHiAT9sjKYFb2o4PA
aKofUCzNLJRZpBpqZPkAogRYY6xVwZYQE4CDO6bk1n3QWGDTas59/IYw3/dtIguLqsodi6pUhZZl
M3T2w+0XiACdOUdxubjbUEMwuIYIEbTjI6IIpW8bFfL71wxq8aDURvyUKvumn4ADwT1PRt8VUI+z
1rO/y7CLk8RIOoUM+r37tlGN0bcBwU3I+A1DqK6NbbC8u3k3lPx0Dq7M5hsqAkItwGDFStYlQJ/f
gKih09k83XKbqh5Dmhz21UnzzS7nHsD9z33bkrni0Ckvooq9sbHobYyv6fnFSsrc5fKaKc2MdsHp
O6i3/GYt5tbKDzr8BpoE/iSDAoAZ1/1iDmjf7S4dd6N6v17T8ZSX4eJ8V9zRLfo9wUcSPCDckHQN
/PtNXe9jhKxNpWqrTGXokviaRyUJbBdynasQoYcj2MINl4PnC8FR1HC2+xyQEnx/oigYoSCU/Hap
Lwj3G9w7WA/TwLwjF3sR82rBytD1vUEW0wP7Zlfrim+oAsKI8WGWfgZU2b7TX2m5IgOkmjBaLG33
5+DgCTx08PKFyW8u92Trfvz+WvYXUAI4gL2j8rj/ldn/oidWavXnvRDcldQE18sSh+MamKGd7wBK
ousg79SQOatlw8ryvHHh8V0I3Kq+ggs6gdgl3r9N1BBtyCcCv/JmuJRSRxTNEzgZrRFWU2gzRWx2
+95HRUfwj4FEhwM/7vf9hBHz2nX1orMu2ciKv6Bov2YKCk3obgpfaGR1BzbKU7w7/nUabZR4NwWN
tmffpICjFkW67x1o8j6OHJGCz8k5wUB9+fUTdGCZEjTKnLMy3EKOzG+vEgVkqcWD00fphyvVav7T
k7yTHR3jkz/ZUHbT/7JwpbCIq5uYgzUePX4jWSfOUOWS00ZxojbPmW1n/vTdGg3NVhTnStksH285
XAmLQHnyBxPFB85gVQXkLjvMTKgUQFHX2WCWuXHUAyYn30hHQv5nJudJAUl8pq2k8lKtsgYCoF0T
Cr8nJTyRZMTf9pXdhWHNk5nmTmyYaSZNM0+gF2oXwNObYcwK0OcoKpZ/W8nOfEXgUCXcahFtCUaS
NuiQ5gCUhS5wbHQ4TtmbsIh0gSVqhQSPZR0bG5aQjV/MAyT3LS8QKQQBYyF1f5hWAGDqpenuRO/F
iLlChCg7cfljKs7TCSbDFBD6T16PKt3phNUoJQXoyruZMiIixZQVSOyurI2nKkXdHsERiba5ReaF
hOdFqnOabw/c+jaLLD5KtxylzmyVCJQ0rJysR7RDpm5QyiurSL2XJeQk1J6CCgQAdQmyKzg7FU1H
vUSllZ9aG31M9MpbU5cFcW34wUKoGkwAAppOghlDYJlbrh31AJS1zTZ5xtCsKxT+Uk9td0xHiSRy
7J7DXFp6InUpGAgNZS3dnA7GMgQRZB1anzSljb3JmvYi+A33zZWDJPjbBajdfDGW9UxZRRaSLbSg
IZpyE03bCmhReFv1Ix7rgW8I8guzyXH0RNAAqBRRxFPg341unv7n327ultLfDwH1/hw9GpTfijrb
oGVVIvy2XPmMHrWQO/q0GXkWy7jxPlE2dhhQ0UcW1D0rS6svBGXC0K5U4IEkdhfN43ynr6ezSzP2
TysG17GEiGhBv6ST5J6ZLHH1JiFAkg3V8Mw6xcZRRIIixZ4MQdT2TiZPshcYy71nA51Rv53xhhds
x9xuo5qLx/g0kX4CzlJipST9ZwAFx8/TPdF49BQUaSsi0rhs65MX4r9pxVXGCyyWMs/kGEpXQf4Q
hgaYgFw13gQiaj3otSE7Eq+cuzjS/H7dkYtkWjiPvFDMT7t5AtrrjHGGDaH8Rn1jO2wlZwJzdgVm
SqiZQ/8indljQB1ILC0hBwdVYp+Rox4PZ6eOjxwyZg6vovkkWnflgcD9SGkUXNg610bZB02dRyK8
olHxZ9lqYI5ajbtutwLGcKPgC+iegm4nTBUHRHbNfyreUByoe+b/EAa6/giZ1wiF3jwxeRUU8aru
5oC3khHjsjcoh6QXa9inzE5f9GJflZPqnv3hwPYrvddBlRu66ww7DxTUe5BlTUs7SZAfcmK+Y5bA
CdvUOO9nHfnjaW4jPlplLBj0+hBWBf6UQTFSaAter3kmT/d9WIdC2D7ys8M36DYcoMpDSH9DmBdM
+ycOo+CW2YAWJnoBYF8vQA8Idd+hW+kAPuhoSivOdaKA+CV4/G1RPETXPQO6ZR0zacE2RFrL+Leb
7kl82HZJNk+B8+y+DeErjMy+CcGUIEmD87ZocKRKvbjZyChgnBp+7nvC4OwB8b4foZKqKjfyLpJm
E+zPgyL8O+MNvhrCdwtP8VVr3RwpI4z6EYw/SiTLi6uYi9qfrzzuYkvtPyfvmCHN/T78CPmFKy/5
BEQ+uBFr85QJupCbfqU9pdHFWvzhNodWh5dHNPsWbNw9olSWjo8qnm5YM3OOdnDVtFK+whXCG5s9
vR94p/H0FHbhoxJCEIS55h0WNWXV60syW04iAibWREbHMzJwPhf77uAdpix58BJiYEXa6sFyLwmR
jMptYQmydzk1aZugs+uZOe1pX8guKJ2iiBzvvmsxiU7IqTj1avePYYLGDY4GyeUQGKcmLMJxJxql
64Lqo8t3xRx4UGNrHEt8cXL8wzlmmt3M+nHJ0HdBVoihTFcj1iUJz3ZZeMJxDxw7OhmBn8zMretp
eih8dbK8slQbz9VuErg/54lcSDXUI+bPwWOzrmee5XstxbQI5G8Q2a0nLWf3T6yWgjrjSfw55u7B
YH1/Swrl9x9XadUR3Oa/cC+CWAugIFi3qHvXHQhLH8hEf2xkgjKm5s4aEne5nYwcO4vimEZ8XHoU
ClmDx7iaZ/NdSvIYcT5LKMMH+N0gQVNW2k8VsooxoGlDbpEWWqMuF6nr16833SCZPkBzNZoyXkhs
DHbzgfcrIjkKQFFt67cbwPZ+tf6iMiFhjpoIuT5PmD7Bp3RYQ3a+21evsZv3L0X3XoSQnxu/tQZb
TvqiAK3JwwS9cdEZVP6LNArGJc6tcJZXvfRbJCNFrMA6MzsTpwLPbmUPgLGfdxanQCwDyhojqZMP
44vHMtNbfwIdiWo/ZJRpAB/iRCXjp9gugAS0azOI3C6JhYaoclhEeahKC0bDroToOafKoPvBaszx
4gC46877U0zpEcwYbIHbvVLhdmJ2FUMf8AIKURTXUYTZ0+LvgezEXlePGZa+x597YEem7c5A/fdX
1uySRq2HeSzLS72v3fXm6sshIiDFfZdIA6AuqU44uLz3bIpAVBKHDNWtzMikjksALW6kli6eKWI+
eciJZVQhB6JQDVwGmiI4eb9ZAeymlotv3VS5lQHL100sztrGEQL9YvChnNsEwhHNSdkwPSi5eCKP
HKoqKshIKHntN84Yx30APDlNnNclnJDv2XYmepnp62Lf9QCICJZTs9MJV9qJUmC3LTB76YdEfNvb
kTFNySLaOKoFTSibYZoCEiVQY/JTLuh4Buh93Nk0OvCG9UvjAVx7kSWmrrUr6eAWE1R/OO4lVGr+
zNYyOglcXx0PTmHjPiYxITp9MJVeK6XM4XqxCfWljSB0FqLmoAgIX5wpFg/GlU5KRjB+I6lczA2K
+5DyTGoZwmlp4PDSUv0QZvCo5Yky288vk6+0Gr1bitdtNbG3LqMfLb4z3itYKGkcp6G4K4H1sZlN
AsCq1k5K8yLAJsGhOL6zLkjizKRghLultjhrPNnyOp8g9X2yqSvYZDCHzi5KWz8tyl4CO3ElLB2q
UBgujbBUdIpntOYcA/2V/vox5D0pCGfzYrw9uGix4DwLJYUbHNuTa0Ar4ISNfGSAZlaEZD9XK0Uc
bQ6itSolE7Vplov5hxW9ADafOFn9+BXeP+hxK2VJNJBVPIB2D0uz1ViiEWN3/xxvNzGyHAw+VhT2
7Qn3y7+fNXqmz3iCGZ47E0ebW3zByd/0OGb01GDpqQoQLZz1q5jkmRXJNjCUhOSfmGA9tg2bmkOc
leMSU7dKeGWHhKyFAwcdeTs2i9hT+SubgTjAo1W4/NZgX7wzPvcgDAZXrkjh6a6YidhyQpqZ0Ycl
ljLz8w/MZxqfuzQyrsyDg8KE1iLSxp1KO7ggvyi7U6lp3O9QyOcCwP8WHWWBzzFtR0gSLlTY5ouk
3PxZEBjSr3jzmKCrv5n7oAzEts3CglavlNZq5Gq6KSsSXZ5VagA9gfRFm1/unUBcQJF5h7Wp+wQD
+n+DOoGWGObXUI7B1LbGH/yBIzrU/Wc5pgsj+pwKSPXjdEdspeuz5X3CC2Th/GrMscdto879uRHQ
8N6OxTTj/Ru5al/LEi96IrQnPCOcaBB++7kVnRjlUkfe6oJdvrCvNsvjfkzkITeOnHfOIabmkz3U
WphwV5UZ11KXvLoliR8rRGpM0Ha4yIJL1D308CvnSTrnkn2uElSzVvlJiCixqJK4jIMxhMdvx9U1
PCFtE8sBNX453NTx9V/UJGI1MUNqPAQhDSRYoqN9/r8EbHOky2l8N1p6WhQJil/hg1omp3gYbyV9
aLsKQqiN+OblzfuJ8nUmcH3SMs8X5vtmBcOMyaBXt3bw5w5ttR9yygTFTbegqSESCR7eM6XF/eGY
VaxMBc66W6Jt7qyp1NYjijdkXBAJrjEAhRrm1YXPU/ZpeSMlFIk0BbsGJYfFJbIbX/WELJDBOY/G
R3tHMHHyJqOKTHR6pYgbuglp+Tuzk5i6MKvEsp9XUsReOyIzwkdZNOU1FqusineBlmPy97VyvLxi
mdZOV9Cwkev2KYxxEogR0zJisVs2IlqEFzWe0YDZByhbm8U4uFnh2Yh2nRE9mkOorRzRg3U4TJfi
szuPoQk+mtHNN+AdKl9sVxYeBH/GiAe0Pkmc85F+f87LsnLouDpfADsdqduUa+z30fM+bMIh5mRG
gVHXiMSUITkr68OTBD1OccOaWItIEfOq7+Ncag++OaPUqSpcsKHoMPkGfcw7mwrKZ01T+mJZGLAP
lNOdcmzaLcpGqUMalEuyM7jWVQ8RZKtd4Xip/cPIDuyqdnBnfroGo0dBmuWQh8tpoSCLFzcw+LCK
mBnzC3wNipjZyBv+to+MnCGIL32D0mHT2kOL8GUvlflPZSZ/Hx3F41EUMiXLj7R9GsVF8aMV77RI
VIi0wFyc7XCwpNzlPOSdaUpaRcKEwQsL10XJeZKBeFDbPa46PWAYteukbIRZU1Ta0+aZmQYBq4Fa
e6kkT0d9P+AI9cspDEkTGCpef8BzN9KcorLCIwrJz5W0qkorUXI92qD6zzJN614cKZvjGtepraXK
rGpW/H4dOjAI7gPwDAnn8Xhwn+YZsDA+P5A8IEGhgp7jovnTMD+RmqwqrRsMM5KvA08Cl4lvb3pm
F/iWqFnky0ieQMX+9Uy+bOwVuaPDDG6dYiAhKHmoYNlG+3me8cbqA5r/Dx3i/mr+bS8CH1HHm4Fh
UzoCvq4YGscmixtCkjpCkvOKdzwEul2q6LzKnNWY4758cEDEK2l/EKfDoELqAbpj9cjNYzXzKoyG
cO1hGDm2TumbAevbOz0hlXPILK9Lv2HgEOCnt09HF8jZLsflz+rLW1+pV+W3s1zDxq1vM0hRUBkB
uZgUK/wRqtIacRDcn3I3BoZN46Qqa9a+UELmvGq7aq9k7px8TUcrAKVbLY5jtSikVKMiOeTEnQAW
1buIXBgHQvTp2Ri3TnUTX7hA+rvh5ofz9A+zpWEjTDlHGykm318eQI68Y5cZAXRhkq89qDd7GhJb
+sdauDiM5EjsFxK5uBu93/ihVCTqEdHxGfN9uwvTLRHSEKqpx7IjNxUlVy1hbFMWbdn4K3BB/28G
b57TaBOaL/ENSQTj0IBnDRyAhenjA7JgHbB+AlzIfEgPKnDkGx5dsQYvZaBvNWH9i/EKKkCNT8Ty
FmnpLBkDjPOEVO6n7wzesaRtT6IrjNq4z6riQxwq4y2/m+0k8s8gR7uOYxQJqK2pVsS+vEQrAOza
Xliv3gHQLclJH0jzQrjsPa+Ds9JEADnzIKhiHwE28i7+jRKJN9VPt6Ds23NooBokVaqesLThAh2m
jGclE9O5jFJolAyRaCH0bTjW+j9WHR7mrKZyNCyDKoxEAD50Pn+vE5uhK+iN3eu0EuaolzI6oZDX
79SovYB8l32C/Gro56d5V8vTbFBD0w9bk9e0Nn1DtCgESWwLHHVIONuH0azPOzefaBqznpmZuKul
tSq7amqRJ8CLX7yGq0U4t002DtiCeNfcxUqOTixOTCOPDsmu6oeqip9zwaEGIvKq7reX17mxrAl1
dQGo8SADRx6b1NvWXO4Emw5KT2mSlRtUDhb6TeGUWn7qH8f7e1f68VLVHWasc5APKT8gf3OjbDbk
BV/YH3o2w5VkJLPbyiNIf04jYmJa4WBvWfMQHv1CpKlx5l2+EGWkGi2cTVQ3i8GpzqQXfj/bjeGD
PGVHLMKmMgSvIrCT9JWj79rKfrpbb3HpY8c9ugSiEWA8/EJCv1FNwAsFDbwrVSQ9ywYv2KXbU39D
ObELx2V//RVxtWk+JzdsrsIxmHF5r8qGAQRASHBxaRpffKJPrkjb5vnd/lAULbkMzsYcrITW7ArX
r46u0BTIlHkzAh1OdqcTwVdipLgxe1Htqkwq9elJOU1+1Pp1NiKFQ43plGx4+LH0tHbMU66HNNa5
rr28B7e8z7NNa7jmWNLABxWIeCGx464IfyBrouetMICvJBX+8cpWURh+ajY9XZfZNs43Aj0Fgq+l
sZn3Hd3Ydw+kcfEB1x6nunnaKXNB/pY8irI3FcngaBMZYAsZw3/1E6IaFpt/MRA0AcjRDmU3w0HU
ha80BoQo8+Y/HWJk2p7j/m61g2l7s1rhTRgdssFOEGijwXflKKjTlWn0UA5sUAhJvS1VLvnt9EAm
9SOgxsejnTH2Y+c0sKvSA8PnSv4lBqKKrPfkffC/xOif0mWm5iOdlJbuySyLqAXE43e6cUEv+sVn
oYTpy0UiUckF2c1721+KjENqMbW+btD5QCZdpZsVVg9JemuSwPpq4XPkQ3nrtTmfVIFP2d9qQ+T/
emG11doGs4k0Or6n1aPhnIbU03krhZaPeHNelYFiluQbAcqRZMQmPO1uSivZJCeowKnM9qeU5hUY
BqpzUMgjcTx15yqCT47f4BAFqQp2xruPpVnUaeULoqNrFNj/Mvq2YtP5E7W9pvtLsRBNdSIgHncv
BoIIjxW+/6lvygibRNXTUHtEp/byg44gIBEZgXqAPN09Y12wC/UeJaIUkyOkyCftjEOivfleKR05
wgNEgQkt++IVyPgpPsFjtTwgq3yRYHswK14HSI1G9p2h/zsz+N6aklX7QOfBeH77u4i8fBnHjwD4
5c0molDzBRdLjP+3hDWyCDsnv7uc4CU7sSBYIG/IlTGvJEi6vtmgv0VNNUR9geY/bMuw1kSNvr6J
UxO4jvE9zXlkz3Hys4vbKqtClZe9DV8K/3Kg/c6txoE21B3IA6HSlgtRGvMt+2Jz38k7nYe742KN
wfRJRd0rdG1TMtDS7fj3CfXsygVEekVWf9VlzX5dAqQEstV0yFFuzFhwJXFm70s+XuEryrDHm8rP
jr+CLBalRE+sLOphd4290cUuyUI1OeL0y/L3GE59QDbuoucL14Zbj+7RyOt16WobjwVNkqclR5eG
tTajQrrGNAugBcSg47ulqhDc8CLpFmVNQsl3Tc+hYygWTwW0xx0MUq6p1xYedWjrfQcceyXIqw9I
5TspyV0GBplQfF9HA1C5vCQJpla5eXVHz/2sXaaTdRXdW+e2MZBLowTOdgNtnsff9mTsU6/9UMGX
bBn1dw9waS4Cb0XKGovW7DvLCjPUJ57293FmGO3OJfn38Jruh9/u2CaawX6yTJq8jhKV2ggQ/L50
FKfVI0UjWm8V6AV8IqrGAYgaweefjZwjVf3piDEcRQDMMw/ThXw+Oc3jLjqiChMLdNTCZiZrO1xP
VhzEOGrHRdJVbcuB7VTZLyKZzRDDsQ2cgN7AQbeAqCsrK2vCDtYNN2RttqaMkDS0yfYOnumOQ4o3
8QkCVK3X/0i6mgWnlhJRhYIBWv74v/+L7fMlhnyqITfaywx3FtBlbfyBoB/n0Ajc3JINUFr52jfd
GG675Vo4qDsZxuTHh3yQNo8+lWLJfcFtFWAVqduadLv3gTtGN/7u0eQZnzg26RhKvAXz5THidp5h
YrzihCvRI83XPlSzsL7EMnSvlXwK59VFauGSssFq3a0G9W65cEhyk6dVJ+kyZPmvKRHuB4/gGT2b
uVbPgg+QuEVyluYWdlMYbfzj+YRExrrX4pioGsyNNAhwE9fQAgCmW061UipYSsSMukngU1aeXiai
0wn1RecG0PLod6NNb8BYkSC5beJRVGOz/vKoaWKis2sbowOCPq19KUE+DokwyESjTtRm+pI0zw2U
+whjzJGodVzELkffguG2AkTN2j7zqbgl7B4PgGjKy3e/WRn4Cvn4BG2oS7A2IlXHt88BOMWRiYd+
+aQDZkegENFJy1Olsbna29yPvCUx7/6YlwNcBh2hmq1LSizDV2u3xZeiqXplBy8BZ+ho1QvffLlL
osdNDG0XuEr5ZOBVSeC5aBl/B89F0+l1sdWWePZkW2XLwX2jee1xmQOwayzB//XTUo+LClcJSuH9
dWso1do14iuF/8jX7J2bdkmyKJr9wWNexuotdTu57gaYPgxmTa4uW1WKib8KuinBpFBXwFWr+vAN
4fJsuDvUl9jWzrI0NNOBkjcygDwPKTzxa/vvtNDaayDvT1hwGQzfaBJZ2hGWtCLyMrFc3ne1pNNJ
lhsv6Uewwadc68LzbopViwVy1E39vJuhTSEBZ0oPVvIgRe6Gu9zRPHOdlyaxI+x+WMmJCbQ4kdGR
HYistj1IlbuQ4apsGBytFRhVo0A4EaVXgxrmcJanh9hQb5FppHf57M8p3AfchbdGfoHUjZm1JP50
3YvDP1MyEhDlvA1XxydrhbUsrKkO3fxFuFHiz36yNSuKXLnS5Q2NFlnKo4S47zYH6kzEghe/+7DE
wPbU5Gkpnqw0OteVlYkzRBr9jSXUhq/R2tVtvX9G0vPoDvQXKRjTgdV+yXptmJJQgmcKMKeD5PT2
deqetc8F16EZywEZF0mID29DN22VsEwprxr3nZvlFSySQm5iM8pvVe+c9OP5JG0ezLq3FxWCKjpn
8ECDrsDceErSjMZnK1ddv+NFBTu5fWSlayL+0ANah06RW541HO18dPS28KkKFqPl+o9doSFJZy0H
oWo97ZniR+ExsZjinWfNkKGRJmat0NuX+EsplW0enQ8L3A7dLl54WlebG0mwmM7mP2UIF7gXWenO
sDDaAyvu6PrZG7m5pXq6VE1BXEls72sSdLtdX5xe3Qtq+Am97S8LvQmQipON1Qz0p28SWmEvgbdk
j7CP6WMPcq6L7LXNlFlrTNMqfNvNdjK3oIyQmR1FHRRuWdkZS3Bwz/w7r7a1itO2hepBrdwzVC9G
Pav3OlnsZ9hZAye/qpELEd3cwH2kifPD0RcufrIMawYk5eAf5QR9r2faGoy+rgrsVAW5rs9kQf+D
/Oqi+aSx8/+fUsCkm6QmLq8WCVYo95HXI06jOvrvQr+BZjcc7x4KJhU6UT1A9HHgO0lm+I0zNezZ
AwePzjzRdz7CIkzhig5zQsxQAwpQMDQr1Pq3PADkzlIx9BypVLSdzrac/uIoi4BZsD5oczIUccz2
9Cb8yPP0pdq6n3tQ2dGhq3N/dXyCNlYEI3xOOcm3mU0YBAVXF1TIZJHmESlRXstQUNqtTuGzcsNq
PkNIaAGr7QLUpHVHFC+DNbombPn8THR/PVoRSaC0ZsV2Ze49XpDg9Fg09idMGTygjUMbzs0ILxjb
VnyLELnQXsTKfBbqlPZVG6bUFrprUOb5vwAuXchacjIezcOLmaPhNtMc6pDt0bbtTLaID9lwMolX
HXuFzHoujKONjrpiwRolxnvlzQL+22Rvh8iglCesIdrOcC4Sa7vyD7Ecb0s8bf2+7OQbz5F4GGk0
waYvl8a+52AJtjAtJhPTJQ2lh37UYIVmku6zeFh/EXN4FME78Iq5saBvxKhkGcYpyZuuOCB8hv52
Mg+XXwiDgRhaAu88cSfAqdlH7rjo2HI7wKdfTS+5XgIF4z17c0Iqlu9xv+DMBdJSQSyF9wdT1BhP
yaqVRLziqsS/F5wdiTAkCbyjA34KvuojPmqfWMrN6XRFplA4zABZMgLiZ2AU+svEqQnFoRRG30Ug
+1oq5LNHbx1coUpeRbVEfv7cIg++O6MwQv6gF6cYRYmOpRnnK//ko/Wb9w/igbU+VcLLgxtH2OT4
HOAMYbG+XnyH5qp8L2P1GVeTGdOxii/ka9syhGTPsWwLGPmcUEVKbjiOH0bcPjcGpgW6y0tuRTRv
zyeBXu4ExT9VzS3K2m+5NnRXOYxGDpD/IvD3n8hvvkhig/+49mpAlilbhIeyrEMLcV6mpEmKLi1p
XIYf2+56tjeL6+AWxMrXXMEDHe3cv0tfqCs0/H1YIojQUAsidEaDLNud6l2ptZv+fksWRgYKyZz+
keJiHqxKqsRr2km9taKKtJF/4yQbDo7APrmm/4idhEZH6LoXrwIvUSiFLa01ftVESmjlo/o6r0uU
ja2YWhpMEvWe32OiRDdKirCu/YHUx78Hp2Tgw3bAMA5q3vSrSrs+ZaojICgq95igWNKzy+JfRkIa
9filYcvLnan/TaSkSAQqkB5rkR1ylBBgMv4I43sbZJacPAbyfajoRsrwG+ChtZgt0vdVAHFtdhEz
WP2KZ5ZumO0JFpS5yxk/SWNknpkyeNSDRUYvHRTcwMfxJWBZDng6pYA9/DvAMbap9sNxPgLnW0G+
5rspgHyU296/fhM7KUD/WFlXOPXKvdq7EhVhcbUj9lAXlLy6M5Er89ERM4tOL9gMESE+SNJ8N+aM
yazLVFaunkjEP1eliwX2tUuH8Q6HdyU6wW2R7r/9zB9lbHz9AbF84XkNEQe1Nlz17v6L4+t8mRwu
+6+OMZOKnHvI/+lQIrNmg5EMVqBGr/UNcKQMGO7yRVcNi579v6yBTIBnyN18dsQzkLcsA7ko2bqp
LziI+F4nJ1h4cjbghACP5aNAojLb7eoa5+rGkNuFvgIs+588DaG9LVx9ggxdZM6HxSzj2WdiFra3
lxcBiraqzyev8KuPp9Y5FnaYxvygwYo9Pz6mUPj8FDU238xQClDB3qY9mMNzpVc2Sg/lh61lrTQy
pOfaRBBFNhUQ0zbYBhpMk6fzdw4I2jH4vHsPhkVgpQAOJjDTfjmy6xI9icv4UGhpwztNDn9/vjqQ
Di55jC2/Cp+gRfyn1DuCwnUFZT2Vtmq3dsgVP/F4MY1MGgHJEAfX5tR/Tv1rOCaHKf2r071KEsXA
ZmTa9qrY3xhpksY/L8MPyjJUOyFl/k8azf02wzSqNGDxfy1wOEucL+XCRxVH/m1CUQfGADGl92QE
LgO2XFWs/ZDO1iC7cB1uxY5eVkcH695of75mNy5NyCy+2AHCFFnyC56qxVBAyXEJKHOkGEu506iX
jIKd9/FQtS5K5bIOzmj52D2dn6iVrJ1RgbdUFDoKwsIUvdqwjOYocCn7A4IoGkvERHY+WZnbcT0D
C20W1q7h3e1zuSgfnmAPI47MbtOd8P6MeppT4WeU5vnk2YhHA/2Cx2u06/vzwGAk/W5KPkGPv73l
sLHN64s9PK+oS80wY966RQsMcTthIE16/vCU3N/QCMxwZ9aVGdHGmv5b8P3FWHLzYG+MLt4JjZ4v
/yDn+mop6hlleOc+kZCpOXIsZOkjNUe7Rm98qMbhj3D3Hr42HkbHSHlRa+Y8aiLkuSpkdYP2lD7o
1zjdD/1Qg9B7IdnOMLSLAK1NbmLPAjgHPTO2NrDRcvIzisewe3AiLNHYuoc5S+ruBpOTAo7IMwlb
DsIOjvOQE0i4c6ThU7Mzxe1tQ0IYwcVZWRamMGJZgXrUWfX2EX0ft3S4HRMqoJqmNg0UDB3XJgCD
nvzBG/w4WLqVq663SpjrMxqOth2uLrFRvztEmTAoXfs3N7xCzAyzeFkZAZrPLVv3984zQzkY7Kqm
urCq9GgnaX7Qj6wjJXK9/xCPaEI6vjFPx9GtWc3N4/zXsecNx0hbFdp8Wl7aFzh6ze8r2o4FQ5Jn
PQuNg87VGu4litABg/Ce2z9IivKyp4qC6PX11hTvQtgNRbFdIwLDP/cx69y7wsDDJmI7EmK0MT5s
q+sGob9qRIOQi96T1lUERg0dYF0FtBYnVAQELj3Ah7PM271P+r35LlIazfQp0Bn+xSXZwx5w48nv
bH+4tX2bkWAYxQEsX545K4HKHiZmajw95m1JG4/ULPWS/qHo2aWzjAFWp9RxscmUmZ5joXgizJQ9
xUV0xyrE4+kePmNRzFQKjkZxu14sprI5L+KOeYF32s5YnjoA9Z+iXkoX0zQ3PAOWtDK+XSsoBwoH
9m33+sH4v0Jox0wzjP42NC73d2hsa9nh3HeHiOaVUNNif2MPYDA2eYuf7e64b25RY8vV4hjD9AGc
uEant7limaiOw8oldIU7aHJjAoL7bSjTsfDHfJ/d/hb0htqiuyRADVA+yqkrpIJ2wRAj/rCb8ilu
/uu6rC+CRHFsYflxHHMZpdZ/sWyiQ5d0V0KN3cCrL5DmdPFBMcfeaCvWpizG3QjVAU4suOyKYWdc
YDBNKmLTuKVYMSFEf9NIF0XiWJQUZdSflTGLX/dGElr/EE0cEYDn0uxBHggY81PtqmUdw16JmANP
yVup+qLYNVZQMf5iZJeb11/72xLWpLmU9ydOcVCukbNWIsTox66SevRVQfgN/EYk68Uk0+Eh0ETe
Ob6pIhz528/GdsbjExkZGwF2uGGOv6dpbxLric29UqB07bmzJgFGEq9BOdnsgDXl1oUDm/uE6+dg
axX+NmZSTVGy4BYF489e2Q2U/1X+SD4p9XLJsH6DpdRS57YBbyOQ2DBRYp2MbkDAnEoXAC7Xqcd7
VPDKSO2EgC10iy0jlQApZoUpMZDQ4siG8hmP/qKI+2TD9tNXRtaae9xqKsWhAHp4xWRoe6LaDo+K
ngZMY3LDLOu6PbQMDy+9UTcB4pStdKGk68dRBvjnSSF49iRGkkVRpc5nWj71lSva5H+fktPPEgfy
7H9kgpUv/KfMc3kei+75jMydU/LynD1X5DdTMjV4yOm40WKYC6XzRzgwaqEMaKegtNlAqO259rrV
dYtPKBKZ0NhsoFRvUUmg9SspzlIsGI2l7PgUW9PeCBhDhqvT9bht+Fgz1lxa1nGGJ/pqA9Sm/u+y
jLZuP9NXLE//JioItdjf/6i0CSBbsqmKcZv8GlKy0+Fwy43Faefnzyl1QlAGBOCppHsasL6M7lWR
WZs5o6KnvOq3TU8a/ycSF44Agok1Kox2tNTkmB/X3aojaKaEbrMRVMem3iAkHYCUu+74oXXqG3fX
7rCdyrAxwvJylrS1ZpKxwzPEk3qjjnbZj6pal8EZ7IDItdkEH7zI0OFVBVDIrwEYdh36ZC3m/mfw
qXYw1qG7Eqpm7oTv/085rmK5BTNM2RwZcsXzTyhW46GyskoYORuHessRQUorRxbrb9oZDBy/l3HN
lKbLcvy9ypGvnyykva01qOJFW/cr+US47yMPWipT2m4jIZfO5TfYx5Il+LdViVcxawN9Q+AYfsNB
T94QZJ9T2z9nzY4atQki5nzmrheQDNMdj3Aq/F0ARe9j4WHnJx4FjioyTAM7uWP0Q9A4sX8GRh/6
9ivKCsG3kWJ2R31jW9rbaM4gmZkBGhgbZviSY0Mwsj/fofco5Nh8yZz8gTv/4Ucne55VuooJrRLX
JJe2ij8GNxlr2f7MHIm/LBB/l7gvJ/B3VONPDDwSKIjhxrSOYuo6cmP/s1Uf6ym1arzuxuAnc6pm
S5Zd27zS3DsLcXD5A1UxPQHEvOtAq5WmouzIwQD5DHAMwkzT+/QELdubex74D+BchPzE9VtPxQR3
W0vaMHLBBNtDo42+9a2JBooR9l8cV1mZHrlpkcAVPsCNLP4Hi4vOKOliVKZ2GTrTyjkATlc7RgRt
efRjkCOwEZhjC7AmNwi7o+xWmoyICDJujSD7T+RqVfVVqlF/I50QVX3X5l99a6freK16IjrJwolV
4N7MxQWhmRUhfx+R/BpUo8Cff0Gl/enrH28wCdDn0d1go8nRUxtKBze+kBK7MafI7UOL6DMqK7I8
QekoxtkZK9sSijMVhYuZb+d5h7dn9v1QfLHMepHP0TkTKVZGAAwtdc6kswwUgDOx9IYIjchslq+C
3rfvsWC2zTt38sy91cmerPfH11UjJX+TlN2+TAokwr8tkXkWgkm/7xe6cKgnfTHtIT6ETp5oPS7p
0xV022JWCnEihQaSe40uPy2zbAhD1p4DBtIkhQ8vB0V2QP6pdH3cG9Uujw1NFxM430OVENldPftz
IdVUAcWdSMGCESwtSFgKFRWjN6AmuXYDPUPS7HKnwIsTD+YWAjeq2yu2hVVxyfmj4rTVJltBZo5k
FQDDeVRVH7S67n+NmnRIuUMaVeDn867q4ztGobKVorodRyCN42mJ96lYq4S3e/QaQyNPvHqsTxyN
BBMQmeutd5a8I+ipwUlNrIXbZ0SoC9TWVLipluhqFzMi+ccSvjhCZp3QN256MU3LacDemRGR177h
d8mAFjtg8YmrT1X5zovqmBjAQ8v8iLMyYYsh5uzRFemZZ4bCJ8NzYnIx1xU2cXfc9OEMVYpXE3st
JFLtPprr+Un5JTU9dLgE+pCh3pdsJhydlLDo5GpkX5yiacQlwhmHc3wkGBPlC5UTCpGcTwGvjoLL
JHwsHFWfwg0uj17d5ICXKOUsE/DH7+N7Zxs8MSzWi3dx4rkSeku3yPFXCbT5Lfasl9OyjeSSzYir
QkODZPatHiuadFI3VzVKCqmx6WEX/qQf/tOzMNPjb7Bvme6pygNAFT7bi2TFYF2VWtIct0CsZrGF
eqzCxUFcp6svHKTsQtDT4ahry09NY3F3TXd/6h+Hta/0RROqgaxabYQKWk91mRvYKvgmOn0UiIvB
Vv8QmL4V3OBSoC7m9y+h+yE04CmQXDS1NWjBX2M+vZd0KHVWtX5hqtj1e3ka0QMCVwHV3Y5d32KY
oltPf6Zy2V88x1qbCuAaY4N58dctj1FIJlpoiaM9M7QpMz2Ym0ZCHOcmYPEFELbUvS0yygbuzQ4C
HkdfWxZ3XguhVetMm1fy2Ufp3/46e0ZcVDADNTTmH/OcRZl3/aHUVapp6o//1vDgTrjz7GHFl4qF
dEXn9eV2wHy6wxV31fiNGnBdiqrGSn69gYs7TWPfVfPCzllRqWslUAqdk+C8n/vuRaW0mCldItGq
kSvIL8YM10P8JtsTjHmBEo4fUJaUy6Z9DHg9/+H0rxoDKQDyXrc9+Ifg3sEmtMeq81UJ+Ef372AY
Oadb14jVjjhsycOIFD7dwLx4KnE2TqlzkDtBmLZ3Z+SmbUIZXLw0Czrtdod9Q/dGZegzI9wBgIxz
0hOTEktbN7BJHEOSnl3Hrn0PFa6okW+32YhX23Gc3bOFqZINicEavbCztLBenWOg+AmoJgGCvT/6
01IZ+lka3NgQyJ5K70/YDHUdXRgFcHWUrDg3SoAIqmrWaZ9YXK2iOL/TCpnPO3uTZ5O96l2/6IhF
kTFXjL3qsH9DzYhJlqdRE0uMFJQE2gx98yRUA0Jt4/TB8BKOhQnmnv2oQdVunAV4dogTccjInNN/
67aIb2F5VeiKPW5Upikbn2l7MokbqjT1oRsH87o5BIRBcGH1lJvSbtX0fxKfcmted7o0voDz+Q8M
w+A526Zz7Hw1gFk1hvRIRKqkazZgpKWABwxhxz5DBbBxgS6vSZxjHrBnCIicwd1FUASB5Zf8r8gb
ehoguAXXvvd8RLl8pwFrlhWhEjEfdxz+FO9YQCfZ2weXBWrFyxGUFyH8BKcakmyF6peh/e+kwS/Z
t9/OmXCrk6fxMFlffSZk/ZpGgWZWhaggkOFeRcbxxa9CZyY1sMNIhL9Kxt3Mx9WHSamj31PJbWqH
aF8mLgm2EcFm1H95imJD/q4vykzUyjjlKJFUkmiwaFFRKtoczfVywoiN/XxN/JxN+yygjcBdZnI4
jtopnI4gSZ7oprqYlntYsSDW3dOZdL//+qzev5YuZPcZteDRkrCLjtlSsuKM+fRA0vORIqTCKRNs
LB+xYZiJSeEUwREMrmUFLV5pOtbSotO8/4wnKURMaRCNcZPqQJCyYR5Q59j7+U7y86XlqX5sPkZs
Bm+JiKUqmOdmKw7KS48CcLWU6eJSfg7AkdmU5TGhW504s4/EKzqi5SNZaeIC4605P6J1Qg7zg4kF
MCP58G8ppd7J40GshRf+qsIefXPXTJQFISTXzBG48b5n3l+zVdeyEF4JyuSH/VVcZKUA3OWT17bg
x2Y6ptdVRAHMEeY6LXfZAHhYSH7gKde+eYA5NvIXaGQgGBIIGG7gTpclkGXw6gqQ1OH3XhIcRqF2
AnzHdDk+TFQlbcBxkzprsMiF9zsniJDbWdACzB2ebUMOSHbc5BG/nQSLDj9duM55JxL9KXg9/mAp
kyXjyUNlYwtUnWHujF0FnYUUx4HJCYbo+dY0FPw1pWu2kuxo8pryuW44rXefe5uIScexl5763TAx
zDd1Rxs3h0GDHC9qCcc/d3UQ/wf+0qty0Kwd6/ridZ6za0tZ1o1QWk+nKZgilCUxXHbtso/bsUhm
bJ6spvxch0ymcMUk0N+4ymJqIUkXZRXduCExR9nKDv46XfeWQ+cZDtFfELP8aQWG7enx2vyVRX6k
a+9t35aVJjXi4tHLT/5Y2/Iavi7riADyVwLo9PbRIeAHBwnbnQDW7BhKBh4g2ZV2goNFhiG0cwSG
MPJ5ndTrfWna4cpEnH5YCjZjJjMY8ANqjbiCqbp+p+oruq5o+7NDlByGlbxPpefhxJcGKINUegZX
qw/asb/JeZnzHzUoknv6vRzSYVZldYY0mDt9cRx+R8F+vWjh6YeOQ7kh9ykaKdlTuCh/ztZMrfYZ
d8tBhYsJ7qokAsdsrvHxzCCgwoFNIn1sMbygp9N/lsM1PeZiPgbo7kWZ5jVWvmhTYbl762KL55xL
NJb10DzWcguqYS7z4G0fyNgFpCspoPCfocVvLvx9M9U0G8pfQ0Psi5NJjxBEC9OAP0j68FThYxOu
Wu6JLtM9+yJN27tnnF3B6ocM8jaghWF3o/uoFk4H/dvnOSAytKQc46rAETVBHvkrCubK2SfhLZux
ZVETlXoqhoo6wvp8wXhb+j5FkypBDh7AvvzN198cAOgAttErBO6ZGLSdgTjbI3GYIbB4YqZ8BxhZ
L2IRV4CNbiUx/aVBWBH/LjS4qYnt1uEI8NvDLQL/VHtyMlWOfzAtQfJBSqm5WreDOSGBOpTrj/LD
4IOERg7Vf9SEhxITXENWDBigr5PzS05MQfFsqgYM9RKT9T/SPtN35s7IxxgyZIUpMI9V09TNLpEK
tuw1DcnOEdqWHfHO5WKPkuZ7GTdYDo1jZvQkrPxQ7vQMgOeM6AT39lkJJsw8wsKujq3n6SSOOBCt
W6QfgKyxuhXeiuifhnllOEZWilQCDQMfWmzi62p4bojidm826csVJ25xe9Dc+310MtLa1lL+XnkX
y2vq5D3FtRqlp3IjojU0Fnc882UA1hXQhqvthI+3tmpG/L7m6zURzdSXgjF86Jar2uHCZYuLzKi1
qRHO64z1zGNxzymb4OscuSJ8rfm2ujLjsQyguegb0lnXmRP5PhPW/0BLiP1JXKF9LzwIbBL6YIrV
shywnjkMmX8fSsDExCTLhPjoIN7jbq5yJbap4sOOCcl8X8wqeoaE9nG+WaHBolejDS+DvuV7RrgV
si6nJsvEUXD+n1VfTl5hfNW2TAESKK98trP+jyX4f1FmX41cLHHy5YTYP6ftNOSXD6eTumDo0IcE
rMuvTyOQgj5Lyi9w3lJFO8QKbNfFagBAnxUGT0rlPwWlB5dDq3Q+RdEwweNB/ropYuB8lQFUztZH
i64VZeiF43EpXRwe6fPAWZtVrhzT58SiEfdeE4m6Bzt5T8gVIQ1JJ6P2cZ2faIWWvoaSWkTcneSK
EgipSNS7lHzgr3a1QlCXOkKMgR1gRmQpE5qtbtGHsF4qveAAFpTX4SoGIOIG2eSfCmEuDp+QoyzL
ZPCE+I3yNwpptliV1bdkpA0hcJWl0LlMzCBoEAPRSCU6rv+x+JtpPRAon+CfoAQ/+Oz1eH0cBdqm
79YJoRx6bmWy64kLUd8VIUfZ9zV5TMZ6srz3Q8nYVVY0b8dsdU/QAPqcR8WIezjEb9IEihcBszN2
KbMMbxLKBSAHphQ47XCwQct+i9rY45Vce9HyYXrUGhC0F43tMhLhg+5SMZwtgHKtuRDfyUkl7yWE
Lsix6kpq35lslTQpx3L2z5fZdexELkNQZ4pMfVhViPhVuW1Ak27DYYQ9DfCkBi7E112C08TSIQX9
u1Ru+GzLOW3N9BGRC+GcGZNDB+UI3iGMfHe1o+JrdFwXFRfey1p4V49TDa+4Y9TGJNhdNvRPLBS2
JaYWGsGmpTILbT/R00hqSmUC50NdvhTyPdLayYtiJESeYsJhMvpVzRFybLzloCT5KKmZwUaGlzZ7
vo5Uxa1xssgptyCU1Y0Xfwh4o3Mz509CKdKE4Wk8YhMEwy9bK5Tt+crAYv/zhDaV9A+BCuHn1cru
YA40qk7fJd2diExCMIULmK6IcBTFeQHIoxWYNltoWu7ETd3g6tDQTGLuszaaVzfqbNpR+Ypf+QsK
uZ5jrYXT7DnZDb3RFhwVeRBKO/tGUXcCLzbeWxG6t3SoYabJtYHynZkTWUiGvWRyBjDrAiGDpPPh
HMJeEzQKSLgVZhONmieObDmBp/HJSAne1kHwNFtTaIkMNfVpftC8131AUCGzHHsa75y+boB/mWjY
iD75yhImp5V40RFK9pw2nuE+8x5SA6faRxVEG+SiD835DC+ub/VQ/md71V4Wu+D+Ds3Dzat7UbUP
EukQSNO3XCFCHP4WPxaN+qb+iwqZTciDNw5HKIWtJlRuhOPIB5Zzql90dEtVuddfqk3FY2TCbV1z
viuQC92CVKkej7A3ySQbmpgKQ4VM0YRL/pc1knaYPlMZJErNi+28OkgZWQ+fqB6ejlGatyPKxEEm
yLe218yS3vlb6NgDSQKhpQ/t9GpDTZrSbG3Yn3ZNTVRyxVhVDuFDcxa0dRd8fXdAuf1CbHwrfreh
/oYw0/zRFSLJcBeMJNAVIJYd7iFo5vAmVwZBRFhtWANucufgOMDk9h9TiK10aVL6vsuNEkMoweb+
0MW+kKw4K37TgNOVqm+oV+kwVx45NWm5pE+jQXuuw/pfaYRuQn1kAdWETrQGgjCOzvTBZ8mIooaB
uHVaE4QEiksF/lKX/7e69YUZN9n5aN0mO4YGEK2ztwUZFiqbhLy7Qq0f0sGHoYtRHWrKscv+0sec
LsdFpOkCWeOGSXdv0hk6/v06iIeSZNXVT7S8M81NivSz8f4ORN2roa4U2MCE+BdElz1qK66usArD
FasFatD03mBgm5G+JSsw+xuii2W3pAR2WefqyCNj8FG6TPmZxSMQLRmL4YgoQDb35yA/+inkkB+R
nDZOYp5yy8KI5J0usrt5LQFk0Z5Pw0X6vqoXw9LR+QcxVpkafSgzInYCkQfnRK2iryTd42V1DPsX
NbvMPKt54B3n3AUT9BIbkx73LjF7J/MOuUcowsOua59OzmpdIlFZqe4a29hCMyXfylrIUWnC3mxi
vk+8vkeME0WRA43EZ5JqOLZa+yTDuu69ytx7dma+ce7v9M5l5RWEskC5/0wlzp1s5Jz+TeHD78fp
kiM33OtKk0GWbdT4XwaoR8d0ry/N8I/XDYAQcINvsN8ysy6LxqkNKX0Z4MAY3mrSmI/SwSpnJPF+
LJkBy/lzAf3lFnMhxWDMdfEHKkBwa+lxjjbZdhJRdhBt0nsJgeyCAO6wF8z2G2VF/teb0UVnfQ+7
rPW7UC9hFw3dKRYDBjjYH7iMpwgFY9ijR7Lo0GalrbOmReR1howtNjMjR7hW6oLV2Zhj4imGZKmT
7d9myxdal3jZUljzilSXvHSPeWx5TVkCI6JxTugEeNkRSxgZ/fvMWVIfRy/yABGvZAoXgV5AygBv
EAEpA1Oi3lQMdEIXLwXF30CtHgup4S6ugTyo3vwMn8KS/RtguYfPnecOv0nW4+QSeP6+N33atjyA
1KFw7LKY2+2YMUThj6QiDjYcTeUCq3qP7tmZLUDtuzDWtMOpXp/8/xpx3MXQfzTOYTHHonhBC2mr
VVBiuAr0rAtC2wWKWjDcqlycP/KM31AHqoO3OOHlNFw1t5J9pV9NuCRYBDUGlXb2LtCGT9X7Qvr8
SU8rSZWhVhsF2aRFX6uxfpMrusBIANQwiM8/242TCmz1Vb2CxFcIAWs2cVzQm2/JTeeTdOLJiXJ1
aMnPNNkfaU1aHiWF5R+whXEtHQocOQdXe3OB8Yyoe3Xdc6WysjXzyqXw8c+WbBxbbdBAk5rBkng5
Jxmy+xyxffK0ZHc5+1LN3dxBnF25fnAcpbfLgdXT/iLOaESgC5WyFslK3TqZpevkLQcLmh32+Zev
IQIdlZQCffIU8Qrccf5NchGtztRlyf/xyjksYqCLHCrrLuhISnqxKueribRrMC0crrrD/dhH0iE/
P1drdGOHN2mweJ2nZT7+thjSH9ZYiAfjS3vMPMH50XgW2W24Z43OiLv9pN+eV3TrlOCfdlNO62q/
JHfB6JMj91op1znvoAkvaVfJJ+nd9Cq6u62ERJXtC6wGkmvhi00sz5rbiP+zEQUMdoiOD2eJzNcK
wOGesv/ZYqZ7Za4u/pKHpOKWYfPY/vTJKzHvi41Pbl2l+/WfMWXrJgXuccw3Rf/HIDohWsHHgiVa
MG4YJMYjcDpTP6eMrEvlDDybOF2VBm3dXG6YSsygry5pTlwukXTHhkf5AbB1DUVZsKdftCC2VIyN
Jfi9mhAlz6pR4y7vfHs38Gl/z5i16eEz9m9E6EA0NmeCk00DjsP2esOiPOTCtc5wB6tDQjtWImJq
ZFb/EKLEZLVE7DULIlE4Hs8sJhZaBcvZkG6x5zXGETx/ra0sJYgU9LBW8dn87CklA+syo9J6Z8EK
kk5t8nS6IS9TSyKnjqYfKB5mJIEdx5cmnJs5gUoER6pHGEkJwTd3161mBA4or+RIOZ4pAJhKVDtL
QXzmYQCQ0uRFoAVbWcIJ0Nf5rJl1MA/LTB0Ksp2Aq9yfX0RV3fHikx8olYKKKyrRgvs/EosaYztg
F63ipj1MXU88FK8MlH4ZcyekcBM2LUJGpVPhS4x1in7CrzlB4J47kbVMICq+aF0fOtSTM2eamSoC
fHQyRkxcVEsMwPfo+qrVPjAvbQELwuU14lEw64XqAFDdjzRIZ8bXSh/i2oVkHr8CX4LOpog9o3x9
LaEczkI46A3c9jgZuZ//6Mtd6o7khlDUd3mHB2j+3k6NEzHVBQpR8RmvGPHXDMr26Q4yDG7UZID2
m8DDOdaZvWuccuWNBWBgdFAqyQ5lfejWEVHvxJrAh1XCVA4ZQR0uJPPhJchzlo7VLNpkRq7V0ddk
bZMsXgP58fJ30rzJ6zhNvsXFo4Xfd/wXGC0jLFUGTypchLQFEIK/xvIqWgH6NquUiEcOv5CcCsTP
O9dC5Nyx5njH200YWqDUxuDrrvHLauj2pHyNc3C0XKwoau+CCEtD6vK/B9AxGmOUPUugacRUjMCJ
wp7OXC+7wptaOixfB5SR8djtZJ0QOWsw9cD7gEL82HSCPobZk0JyYA1d5s7izp4oSbxvj2kstH6k
NRMiOa3yTUfQtxN1pHY+Pz3yYhzvOGxGh2ETXzONK3jnsyWojuWrHjLfr7BsaFoRo5UuppLmk0y1
xLLJb9JLs3qNf4HI2dwIqy18i3JKfivjV7D3wyPdrgiO8XPbECuM0uYJduScz6MhBWo0rM0cYndS
I8zWdZjG4+VKDQb/JsyYN0cVeF5ozUfbEAIilw7QXKMZf7U/p1kenEDlE7YegIS1YwQrBwzJEh4F
zkI8JEVJVnbbZxIiG4LIiS2/BTzHSzodW9ghWYxOZHX2/GuAOqwHPZh3oKVSAc2s7fIqSPl4sgig
pNOl5JIj5sJQCSJNOrPyUblXsOZOx09yZNl+8+aqkEMIj2v4PLkA5FMxoh4UVmO7YddcNszHOpTw
pLumXSjJi+6DVmSxISRv1QEkmb8swn2YRElinZwMI8KrPRJkEtd4P89+7XPGpkWQrLohz6/Q6IwU
U0PfvI0skz1z7FJRehJFIjr9+dV9sblox0ulNj7NfWSIO5vS1+wUWfErob3Etf6pi/nN7BOHHAqK
xepnET7rHwSNwUbhEgB4S1Qo/s4EPwiSLHVwrlchwa2G7LqqCuid9dNr50ME1shXRgfPQgdqLbpQ
In3imo6ZPBqYvr7taHFA1tEQJfnLPxB42+SSYhF7F6bVuY5/6rB9+z+B8HJ4NKtY+feX9l1ioGWV
oAO/DNsRy0EqnStZkPqa149m0QlU5Fah2CXaSTzi3Xq6jREkacLbRkb6JHOP3TKj0Y4CmSSqKKvr
8K+ermAzM87+ealaUTPDdVjxZ7lOmmPb1ev2hw6A3JGsVT5A5tfSPnIYeHejLRVCw0JR1Yo7iohO
NTL1hDpbEm7q7rUo3ZeFwRnMeLjVxSo9oKIVUn8VRGhAtjRu/R0vu2MWyA/srEyl30m7rmL7WFBN
a+wIspU3FEWwxMK6P2Ivh7WCO+IopzAspqugUq+0graz4euLL7U/2feKnH3A40Igtqg2uQHBWkbj
y+CmfEmceYCD8JUZ/Jq2L2CuUdafgJbAh/7jgtOG938nu3FEEQpIJFT41MSPimRVi9kX9ENehKC3
JF4V/NWm5mdt03POnLGPRlgKi1Wjd6MKEVP3PHiw/YbuTcbvkdFlbKa5bHWnaMifjRJNf9FrS1Ix
/zxLTUVAYiK1amBc7YTsDoZKImytiwCoD32/6cqUMSjYcqDWRmSXOPUCyj80vf2gAXqH07IIYKDI
HNslUYx0rQmQXGfqERRJuiaRtC+QnknblnvQdk7anzoirXi93VwjXa9pHFrikyUFz2jyN9bKrmvY
gP13+fhCquvadi+eQKl+a5KWi8vt2PrBQP1cNuTjBk7FhclLI3KOUAf/EjxAF87XhhcdhajcpuDv
nvCRzN4zPB8NdXakqphu6IyaTzrri4ffCe7R4tHdH/QNwYDD/UE09i2j/BBjN6LLQ6kmVF3sBsEu
ifRNtdbKY2P0VMAE0sANykC6baQqHfQ2TG5k8GPat8q1lFIK0b7Hwf/1OpChz0LnCV1j4//CQ5s3
s9joiV8Q9vPsJR05jNGo7roLfy/z6kT+ehxKiTdVb2qEakYMauAMQTXBEAhvw4W+P4C2+2I2Ixh7
cRBsXbvLopD5VTA8xnlDzVBfA2EU/0XiLDd/YUT0sjufiCj4MNPgXDTsVo1RHR+CD8STHvoe5cRo
LkdwUedVJuIyOIt6tPHOEjxbhnqTcw061jVZmfo5x2w+0i+R0d/qsjWnAgt+MD2T9vTZh/tlXxJI
nstvXKI+thr2ZMCe8dxFCDY7GLB/9DwA8GcRRY6fe3GwrUT7CBkmofNiycRU0a9iN/eR8LONMWht
KQjnZkMfTbzYq/svgoZiJaF2bIBe8TqSYbPL89WE6eIhAqzw5hnw/XaULPq7FvlldPFEok75y8jd
cbHQY2ojZx7UX//HV+VWkMdGCPz9LoGQ/dguk/bzvARLbRb3oQPyXacOTU1rJOHZQi7GN2PGxRb8
0nAgdU+NT7elSwRSsEn4zqWJxPG/YrJd0SNhRJoBCqQKJ77wY2LTW2eBt1/qFmThRAq7+ib4crPL
BIaXrK/MBXqkSTF/91JfkY+ShMo7wraLoOIj1v/fsgwFy30zjH9AWZTkpoestsUyp7JE6qZ09BaB
vhek1vjma/deXxkcouiePFGB3zVBeO8n0eloyylbnjcm6xFCqEmcMKmzxxSKvzZ20N83SUAq8wxC
w9i3SBGAK9GNtjJTMp73vHcsozuX4GPX38SgKJ02FO1hj0HsavLMuoi9TtxM6dc1FYrEhrHeADDJ
xzM/pBYMc2mIS8J8G+71dsq0QRpwUam+wtb2s/woS/abmhSyGvrMGU5eEWAzLGTlNeugo62OsfIU
H/sW86lhTKElbzPW/5nZJLKxYwm3I1Q3WkXWSpbzhxm+gB973PtE/cim7LvT/YTM5iqCfFUn//cD
928PRAizr5gygNpkhGqxD+HaHWm9DPl8HZyBOZAYacEmnSmVFQ3SfBN9FTjUnGWHfdPFDC5gCpC5
z3qbclmTafaAeuH+9DE9Bd8Si6V2NfLAxUZhTFErMypGmdZzdOYnLDCxssuRszekWDgTmaBljvHn
w/E+EHgvfUeUW6FAmP32zrHArbUrt0WZngc71Qp4qc67EIWoaKz+Q2McIIn3n8+q5TsnlxNx5x7x
kFmyb7kGUwNKoOArdLyfvPr88AtnIPDoBQgZDasPLNU8YQD6sr3rw4XtDnO+IAwx5KZdT4DhApvp
wwxgkbvNKy75w1pIZ9YJ1b77gJgp7UZETSEU9iMRKxPCrnfqhv3/bxanh677Fmw4n9KgqNcVdtXd
1AbdSA79VTHJNM9yOHDvhrt9a5nUV9HXZzh7kCB1C4rlLDDt2S8dBRFd5JVPj1/OkIE7Nta6HxUa
BDFap8fwA9k2lwY3I7kPcYSVq7vYpwveZXSKJXM5RRyH2LQXBb1u1aSirlEhUQS6W8O8B2o51xNP
31BuQJTzXwowXKwfNJPO0yGJpN7LkkeW1ztp0b3znPSkNiI0kV/TCPDqYKASGT+wzPm2AkzIFMOi
7n0GcdrZdBuFEhC63tuM1ujvllKYqpIsoNVUAL3yWcSz0zzUuwoflK4P0gsRxB+Xbs6cv3Rdobae
Ry2z3U2ZKnbek5WINWxSws3FOnlN+ZouHBRms7Uc9TmXNyaEFx37CZPiViO9pTLkML35s2Ndo4qr
8Y9rbgkRNBrQ4GgqxN65BGS9A+noDBGkd22i8dHpMtrrYLIQxNPKkqp1uFnx5bFn+ww+HOpQCQNC
0dlJRJYEcFVRgK6T/IGHC2xYZpXrXDXkVOfEW2QnqdN6AoQ8TQvyHgiNIQ8U9Xfz0bdhDWAZSwZB
Qhfp2x3zg5s2YIcB2ZfkkwF3K+vX+o3NMP2zog0zD9AhRV0d05L2c0NQKPrnLQ99ah2y5itpEwG9
FI61U4fHO0I/ROHjlBwLy2TnCWIA0AGq0wFGxlUH6GNHcLCRwbnJnDrAIZqg/uLR98+y/8+dj4fX
zAXVNhZ4PhAuz4Uiib2kXR+yx5SLlqUuQCEpGR7Kt6oxl4AKBbi3tyOUWv9Np2RTd2fb/VsYvoqG
ZK+u3d7Eq39ngkXkWkHiFfJsKxSBAslFBG5eBjIQVgNIb5R2hBhhfInRPiTdJIFA2smF+hEygTsu
En/sashWZ7G+gdc6JyU+o0aqw7x3o3QNLdFKyCBAXVj9faRBytPwzW7NgAFY5rRQ37HShceL9ceN
RvT7jaWwFl/V72/filH5R+X6ydK2iRFCgz+5ot3pkrDgTgPsvewfsC5beSjKKMgvm8ryLJPD8nma
80297RqNRag7X/Vgo43y/L39yIRgivaoVQ2zLxNbq+vfo7tyhUIyKdswOeaVPSIiK1ivJ9gU6YTR
GRLYCyR+Lz0TJxAfRBkywRvhb8HXPGcXM72PPdTvA3gy6wajLcnugJGBoFrjJfwrX4IomrB5yzxt
oll8KnPljZxJoRcEnHdE7/dRFKzjD4/trb3PTw3YSJKp726ZK7qVf2BtX1ZCf1m+96ZC3wB20Kf0
Yg1NfPW2BWk9Viq3DZmi5WXh9ToY+bEhZw3s7BEbS29IYG0CZvOQmUe2AnH7jqvCpubG/Koac/OP
t0CX3xQKZX0MYaET2Weim6q07HKNWsMMFLgUBxRQTrNkbIqo85N6dzc/f/6Tpf9vgqIaZ3RHntwH
4zaY6v7RTVYzOjAdzcSHeSHUA5wVfQywEWRG2u8H32OLsjLOPOcqxJM2KMFFEUsTj+Tc+4FAbiPX
+r5I7qWP4BKUnQ6qiPj2W6N/DWtp2sgMs2ZHyKWZR+w95jHmHZCAO/8PGN2Gaq5B5iu/saaI+W28
SkE2DdtU8mf72VQ38tpkkyii+kFT6ly4fzh7kuoyWEgYD7mJGgf60iMINGjn9QiM2Rqq4si+Q+ZP
A/X3zL8ERPuJc6lrpeaFZa5bl1Wpv967+qt2R5ZbhWmu0Kti6yqpxRAh7FayOmoLdle9yMxVkoIt
r02u7JW4E+TXoIawBupgQf3ZypjAqh/KRFFzyz3Hna+WdWYJ+fpKoA7yeRTaORko42g2KOvqA+Ex
U4I425ilaAxEiWJW9KHB/vaUh/lpuQeD7I9FXBqhooTTwIs+zVAcmtArH/60eaiFMl469EtSoKKF
AKOFUVtOhpGBXq86/GqOvE30AQi+ruybLXQkTFHKts6BeA2F8T0XOxRk5z6w8nADCxmLdoC1Fal0
1Xx/ACuOOP2GDI/3B63kFE/XSrt3lVhz2lK7z/NISkoHBS/mGGe3h1pTs7ajrQQi9jXmP/xspG8Z
QWFe9TVid+YwQOcJhL3KxGHF5qigTAOwYoMJi79TA6ZQHgFzD9eihWOys4JjjQXFbU4Uic/xHn8C
saDBWd18L/mmfsisUQKi2NBspkPJhf6G2XBzS7n1NjoBqX8vJQuhozXV0sgC2gCl5cgI08Qer49h
Gwg0VWSzzhSpZMptD3fT5AGfIbVTia5yEKxki8REzWog6Zc6p/T2pDtdHWtkaTQmxJ3G6AkXJ107
6R8uByMgmtecHiMG5hxC2jOFe18aGj3JOgS22BcE1z5z3hWG1jNcN/O/4qT4Jt2s6mvVJzg7mNhW
BMFzVkSCrxfb6uUWhflwm+kaUPJpxjPysJFhE8O8sMeo8uciEjqFxLqgefJywP/ythn8vWTrTDAR
sGbRGISyacNSW4yPgoywrddSlBdn7swvEhWmIeGHPhlgJq55S6nZuwaABoX55aUeTWjOeZqD9exC
OSCPeZyAf7uVYsHbzAatcRSwIWMxMSqKQ6eDZcViiR/0QQ6b8ERlnmNtpoQcHyyo7492o7OkrTCT
aAzOxVv0pRGk2ifFhosskBhWtvS5aTgT1j5TKTOVn1slsFOCk+OtBUwOuDyHRNNxd68n0GH6DIUn
D+ydcAl9YPQGCGuGEqM/FQzbgsQtosdRkAlGEvQjVs2xfWSaX/Ze5Ybq1PB3zvhdnLuWPQ80dEPs
Q+EDV/ky05ZSv1HnBi19/yFEHRWBTc5MegbIi4kQfiGQT07sOCrcsnk6EDFSrhrv5ImBlLruUGFQ
teYzSuUvbNZRV7qqF72ijazBFD6u1VB2wfOrzV7nPhmLsbEulwEh9yLIgX5zq3fQKVNndZetA9c2
dIO8CfxQyFnQgmooTltb4BR9uUphaSPYFV/QmpKAcNRPpSAOS3YMCkhqqV5uzxk7ZRSAg/YGJjAP
71I5vO2/+Oefbtf+8YSnk0l0skDr3uOiku6JahdWTFjqGbebbsgLzXjjKPsHt4WkJKlcw1XZwDWL
0zouSTJAMctsK1PRm1tjGtUNc7ChAl4z99YGIkd+upes1MAkTU0RxHGJBA6J3vuwh2DWnyEVqDPa
EB8rjbXGA5F9yFG0GSJeigJzKzbQg/dknsLkWh3fGtFccqWol1EMrhk++pdLd/eam7QKULHA8Dqk
BTp3AYLHdq5Ctfmpe8WaxmK+ohQSHDSGjQO6sUigjnxEMqe9wETuq2pV9v1IK9tBCaieRQmANpUk
UMbhgzR9jIDXvINx5s4zaKksH++McC7eMyf5kwCgYJ120UE0GVnGSjs1HJh0Oe6CUeo1pKqGqUsn
y/RT/cO4arn3wOKoPdLc3zjdPErtWxWfVPk4bKVs/Digc/9F8lLw5akFkkI62jfzCnnY5S67+TSt
7A5NZGI3lOURjk4eItHWu0gQP5fzPkG9y77fMfhf3jK1zDrYdHJ78EykSvlM95D7o5w4C6cvDxDu
RenHAoGw/TcLBNsXJQ4OVeRmyeaVwGzPrUU4gpUjXPuWNXZeZr4U3XkbOtQvfwfvTglNtgga5uHx
FCcMi049hcnDGVAXQ/ZzuOJn5icCl8Zkmgghup789VkgHrifzxO84Q++SWkyafoLKoT5/bxLxlTo
k1MfMC83iUpzhD+4N3olzPGjVXvmBl/or5Wv3A0O7DfwQFbZb2+XShyt5nmG/sLSUaOWiDdjUuSj
5zXtvQ7psxSQagOE8s4qFsgVal3w7q1wE/YbxcTYdKl3RKBu8QJjn8mezlHsbbRBuftCY6E4w2l8
b5GoVMyG4ZCu6hap4pPE/HWLOBYGr5uhLeCa59GVotRHFalPzFADELSBmRNj33HB1BRZl0+i9VD8
Z3kJO7vxnUjJYWX/GWmLews/aQXf6FfIMiY0bYuMdKkwxxtkDg4MlPBPhttogw4YVE0sjI+IiV+7
SHg2WsDdBbkbyGDLh5gFImwaPRXlgZ0pRDjdKyoyFGu0pG+4ylrd25KR42GmyE78pUtm7wSkcf9n
ZPvGEMei9R/RNgzFfSbfW8wgVuUpGxFhGC0n7lAQqT6XB3N1FkJ/lV/farVrfxjI67s0zR9SonT6
7GVeknqx/MS/bVlHYct0xZNpBDTPxxxK3RVNtzjb3kEH4Y89XZnq2UbiyAEok14edxvNf58oeG6e
nC7rc6xwnX7bXIPqWwlKifWrUZServ6bpKYCfid6fOn4pCFc19uEIAWvoSSsTpuYwEL2SN5BElUw
L8hBc9Y2CxTXwusU7Pu3xBsxgTwuD2k46FuQZLy3xAztxYaSCS+UiV03Cx+muF1F8BDW62TO8Mxc
r1CRh5+1NnnwQISv3+P4CXnyL4MCpCDYw4CGOUcfxnCblQGZTy5pl5rWT92foEvrIGNB2GIcESbU
+ZD+chsKG4RRDaGsJNIFKhh7o3iVTQL0Gi+HxNh6ICBDQ6qtFkwUmRaQeKF4c3Zj9OBHS8QiHI08
Of4XCCrbR1H4Y8E0kvNM5eBTP7kOV/Uctk4quE/lUOc+rfejt79XYoay/9h0Pj1CSdu5/IjZHqI3
5p1GVKei5E+pJPFZDgUnNHB1e7MYP45RJAyj7NVnhZElptGe+nPRkaEeicfiToAkfrxPs99ts2ON
QztatpI0aqELDn3JqaR7MVPJw9EpJ0ZeEVbzMR/0xRHbVRv/FBtNESFu0CoIsDeQQrFBDO/OevkC
zrDKDh1g8PcSn6Pwta6T7Q043yHjQV5PM6iSjJhpp0lE3M8uV5qkPDySJ+BEDz5mX7yNqTwTLEHb
V00lXbctva58vqZQsp8HetDUvE0WKmu9O9yWroNsWPiXpcQzIsVt3syTFQ1pS3tne1JGUY87Ko4W
vc/By+VTpRIgmC6nXfxW80rUVYBWGYvdUhEyuTtYV/9pZf9fDdQzYlGEW14wZ0jh+MCnX3jUgwe8
S6O54E6OrdzGgOScm0SwBkN+Px+7L1jBCZExyA/yKrztr/91JMlog5xvpJ9AqDjJtlYPUQnEFLDg
MZHjvgh7rT+CE66d8AkY4M889Q2/MKAK9WRGOfa/PzUdTn+ffy1pPprEoDVenAE1lrZrgjSTLMX9
jjvqpE4UbLs1qfeos9Urqgq8ApMybMJxY5kvT4Y+leSKTKShVyeRoU9kCR5hovnmmLQ7TnLzNidI
1APFWQyB0hOxoEpGwxY8idnjn+N2bp+OMblMxG3MmpRoSb5WsYC9JDd0vEv8CEnc+Eix0jqLMmX+
BqNNgjAK3GdyMaa6xXIUtRjSjyi7P7uo1C49Wp4JVVbWWw37JHs5biO3SLbhx1OmV/bYR+93fSb5
Yi6+zYu3DGJxluguMWCKiNO45Oq5Qu56fjUMGtbYSoHyaICNgefpLqKnp/UqEWlH82qSFv8d/FIB
+m2KvKhsWz/RTLRG7c11UD5SKNvwVZQG6+UBu4VPbMJXGu0ZLGmSzc1tTC7UPCO/MfpHGy1nC1Wh
sfwRiGG5DE/pwZgP+LGi4OtjqfXeQ09R7Dmo5agfgOp/4k1fB9hztisqx4YZvVwyN+tedPOrQ+ou
uFC5QyD35qSRuDli1Dpye5FD7WAYPrhP26SsmgAkpbA5g3ibcVPj1tslTOzceZjN/t6wueXZqfUn
GFqcm5NgXgMK41PVfAhdVzcZ5vHGDSGBcTMfXd1iZNMlbPJ00K72gsJrvG/0JlSBbyMv60WGHvDb
mfLrSYoiav4bypWpyOvdX3CpoaUEWNZkP9hJ1mseNed1vybchZSqyWt/EmpX+beEMtQpdSHebaN1
AZjzfr07X4U04c6sTGrULVwAp0wZAmkAT08XA9jFg8TrdFzf9Ou7KJmUM3M+qh2F8YxpJzcHIyas
ub1xiJdV0FWILXk55m6WWXjPfOn2ksDh/DmR8JR67C5HDu2ou77lAH9R+Ul3GjQxTPMjQQxEV8Kq
cT6/gEG6TzpaHPm0Yo5RexRiWlHrglzRjHySeZAG9y3igkiJsRJVCGrVt9l+5CFuwA7y7OXt7uYt
GXe3rcO/dE49eW0jJN4QS/qKmyCu2dGyMiJGCbr6dVMu0p3ciOo/OReAKniMxHtog2WVnVmOxFXw
Gq4cMD8AtirQdq+d6v9SbmoRi+rhr0GNjDsiC1/Tnzzv16POgNREEAIksV0RSRJhDCv50WYudtVt
b6qgXVzOuF6eFJqetNCM/lWIrXiQWSYMJteZ/a7Obnf3rbzg3wG+jRS9SGXI7gj/7ZnxlH0sdKpj
IWvJPye0EL16O+dTlWVkXUsJ9mygQ6tyHXSej/UA/MrjUuzFeVDspESp4V2oe9TaLcbNmvlpEmQV
fv3UpSOl+DMV4qSp5lKcvaweYgtjv2RJ9deUqC5iGJe8j/Vv3y41iuJGonCMcGmianOz7sunUzco
r4nYu7bmYRcPwIcPtdkCO5xX2p3lW7u4ukwPrQPN4LEQ+kIOKVibRusVcZLGUtf7S1lBwJe+IBGX
xFB41mi7gE6UW2FLmn/B7jCphZ9EwHsN4W5xd+92lNbeCyHFz2MrcVlEr6wKDMm9hHETXhlvO8ns
gcDPctqp0EaEWUf7aykEwms/XvsXXe4qC2dRtxX2jtan2FJY4jQoCQhkOoITbIqa6Six1I1l6RMt
KH+KojltcsaMytCa43XagD9vab81EMqEu2XUfEpsfcSMF4Xd/htkD3+xbcFJC7ajqnmoXg8ifClz
WBZSTVmHoCvu6/3WHU9gpITGqYY7y9fdFGFSsN6L/2VTs3uGMr6HaWsLBujq69b1AAly/Yy2GFOp
eoFt/3HMFe81+FSsIWWNxWFYglvQ1C2d3N6HeKH5hrYcUr/1znD7CUvNpdNUVpZJzRuIa1F+tgbg
5qJbbGdNdQ1iY0hZFXWsMOEIe/UgraaoRkKSoYRcQxqEzzmYJg9UojPQRit8PUuE56EMNtrPt+h9
wrNKVgU43GfuuRXJicd6RzcwLh1/tP3EcdD6MKp3aPR6CT+ANoTOnb65fiCw31sXmiVN8/fDg5Nw
zZnhgWv4ECJFjrXS1r11ZYhbNa6FZpUt7ZSbkI/ldUqVl+Q6iQK7sS8G3C7IAd+v1dAxPkdIi4i+
5xeKf2qlJ2wtp/NP5h/x5/FW8nOf1WAI9/eP9t3dxoUhVr9V2ztSmrR3Vz9/Jf/owC/f6RUMBLZY
Zsn5rD59/tVnGXYxAGfIz05cTowe1AeY3rwM97cF5wafj1Zg0PHPkfGP5f6VGJVn4nqhm9fNpAmA
8PV3yq97kBnrghxAfupzdF5YLXoyfF7fBwR+v1/9xCh1vF7CA6KL73p1iFvy07Fmrg7E6uNXKna5
FuYdudvP7JrQFKoESuFl5n8VrMZkxbSAK/3Iz0lGcByPOuh9QWlVH6VBOWQpFnFOUScoV7l+2gk5
H+98YkzoOTWeF27ja9xNEZhhHeBNlqSNZ/cGSytYNlZgEapvJAmy2/38VTnaL21CtFs4EhR9ybjV
dEM2qIzKjhum/p/lZkdr3NrufWY2Bl5uw/M/HS3/DCrS0zhZXaH2RYvad9PBnaogqyiS1XdgH/K/
mWQ7ou1ctFwjpAvdkqokH6Yx2AZcnFpqYwN1MM0HWRnwrAy9Bxmwjll+StUxByGQw7KWFlNLDYg6
ptIDp3EALg65ls6isNC56HVSUGxUzGUY5zAFX0g0fu/YBSe0eZ7j1ZDse8hFTIVsgzXA8lbzrf1K
S8bGxJCmp3X4Z2ocqtxGPyx+EQuRirAnguPDJJh1a/hmk95vu41LGAyXOKPbRfMUxs8bdcjCJTeC
k2tnUFJfnrKWV/6qHGTlxjcGXdeeSUsjudlp6eKaZ87THKTH7v5KlwA43EK97PnwqGAxaoWjBvVD
xB6pItOTm0MECL0Pz6wJb+V8DWCXJyETESLgdQb1ucvPWbRtp8/+cmvJigo10sZ2HtfhEkahtWp8
EpZil4QcqEOmjh6gwzmo1jyf97Ni/6mugeN4bMCbb2IVI1l6uwRUG34C+dyLbeql+hz1cQArIWQO
qxd6aRta30COhusp2n3w/ppynQ0C+CMZbHJHDKUiVRRyLULsdt2Y5Bede3I8JIwI3J7Ki0gPu0p+
KQzx57Es3WFh4vM+U2W0yEXNzyT+IXkr+uX7jmT3+9f6xCn11EyndvhuGyji+DfecZx9/bX899I/
4K+kAxF4QQzX1zOrDxolcqG399i55JOd5GlKI7MIz5iVFaU/NlSO8ApxyHQRcLlPgLIqlayDGBBW
vJiE0GNXoS4z+VS0fqwIVq7l2Px0o5zpEbfOVF+Nq3XfQo++uQCGbLEX+XOsaI9KoNrIWTpysIfZ
TPW4gAseHMJr05J6F1iBtus7D827Pbivr3bZK5J3CuQeIDG2N+AtvrUDYTlAik8bBQUdPxPOEgUt
XCVebPLbg2k+GQ+N8cqC54gXV7/TXZQi/mA30g9uBZTuzsSOjjqRcse0rVayM57BP68+iTvkAVyz
P/CQaLXzjoah0rG8OG2Ix3hUhMXJuEZeMlycA29983LG7kTlnfCJ87lXM03XlvAcoE8jDS23QktH
J/0N3IhqwFdIfj3EvbFQKrBczkbqWPaqvOqAR7d1yGF34VrmO1vMy/nRqi2U8zYlGFFsbJVXv2rL
LzVseq77Z1tMEmFWolNf7O0gKJiwFk6tn9d1i9KepjBU70sjrKyOrGBHf0fPDXmJChnEuMZiSpWl
vP5HnuLVePIxMGrd2dMGxe/pslMWSJ7Y1gx/6fZOiamOhE32pezO+t33WSy2fi0mvd1bEntcItBJ
U/5vvp/IFotKMVqz5KtcAkS/k0PWh3aPG82438r1qQVs9zZi0qRjvz5fnGS4OoRQ6lN1nKBkxm1G
aq++D+nnQB9rh4nSl3Q2I+A9a29LVVF/0URVU0plhWcdRtAFRjbbMYu0dVLpedo4Nbnd5tNqiwcp
xPhvusqmSTkDhZxohIFhS6LmYdrc/kWeOlwMfbzpBgLnk7RTVIHIF0mPKN/7ESDChE77ppHSfARL
XBA7jzCSBZ8m+dPEdWSfPRCVI5Cj/YGKokN42V5qff26pi6s9zkKKLz929Grr4CAoWr147q7ErDs
zPL9kFBBMJ6I0FmdZMEeyawiVha00v0OKD3lAUtRxZF8U//mKBJJKhBG55skhKf8CiWZ0KKV/kuA
ml6FAIHj7bI3vAIyZ89zDNo4JFTBuVpEAdlNiDELjYx94GBJS9sWOY6Rmpuo/YW8qoG/6iid6TTC
lMZda6l47U8MwzZ6AEWgA1Mv5h9GdMFDeE6demo7hIn8iNtTrKx/LR4aJf62gVsyogOVFZxj6f8H
U4fkGkqy51bEOHuO1HAHFpjtHJbr64OcpydAe2PT8szi1DB1xH95C4eSeg8WIAcm5JvzOa5OMU3A
BuSwrd2/nAMjNMNfWN7NF7aqPve9d3i4a9BNKcH33miQve8UyCVj/1JIgcg/o5ZP5Sndtm6rSoMu
qiQiJxu1SeviWbxrPsye6deNjVqCV5NGH9TnEDdyHRklc0ouDeHSYuC3XXAr2Yt/hwxThVd72O1K
+FCQY1QdxMCa6p7RSOHDws/M6anVqpEa3YFMq2FbSQJY66/yPiQji19beleKnboHWl/xRAUcPAbL
GGLXzZz8mx6XINGUOm0YR49gCa7WRYLSzHBzKUAV4ObqDXbYyo68vFQQC0GLhr22wBuyWY8S5TO5
uigZC/yFJUpHgre9CbB5J5nyUmFKtJvZvGdHQXIygNfARbA/AJYTdy63X/ceiHVxLELIos2sK83G
jvdCyONqMserywrQIUsY7ABCWN2HKbs0OstrI/GjWcCuoULdK85DQwHHSS7ZH4qH62Blydgk4ziS
hbD4sdOmB/dRRP3yiTRzQHH7GnrzvmMwgpuwx4IDt6Lge9pvPwI7fLUe/7WhZCnW9OJHt8N5lR2T
NSCb13uDVxsj6iiUJEPO8+6MgrSun823eaTXjNLOK7vncaY0OGz6ApCKAHShO6tJh07CT5g7Pa9q
jmK+G+JTJSd/rOOUFaRS0bcNiQvr2jv7dKeoangPyAynEtK4+jM2mkUtVjz/RLeRE/ri1Q8TC/Pn
q5dNRL17XhdsLOerpSQJ/+Xa4FOlPh8lep5oxIvSj/F5g43ctR9OZ2MPV/PhyeZrwBBUUDel0vGP
3FEQ7ZtJqhNIvFFyppTQWuyB8M5X02f2s5SzTgM2noqg19MXlE8nv4URA01T1uLLZNz0s9iOFLDJ
omXKcMWCQa/ZY8YoSQ74bI7gDLSqbWnruW6729ijNmVnsbLA4b8fkVETpb+b+IeuhVnmPwZ4cGPP
VHU9khq64t8/rGhbI+f58e9TLVP+gWrpuXepUKsazigN0WpEogI6bcFOdd1jmKaQeTppzks41Yhv
umXdHLlzERNIV+GRrukIC2FzQ8k8hysplwFlGz2Vo8F3YZ6I+2PTlNs5kfNHY2gKzGAUNvH0OOI0
Zmea7VLrMYUk2skl15V+XlatWlbmn/4QO+bGksQSIuuuZA9QZ1MLvism39Gv5lPr/PIywa4qWSIE
ybhFUShEX2/ndFI/cR3rF6cZoHZgpw4v7RngqRPlpCtCWAQaCA7YUgmY6AQ6SjllXqWrOJfJxkAw
DL1+94Al5rAl/EPK0N0LhnaC19uQecdlhiFJC2PAFIWcCywWME0YoMtx0T9Z9BFMkDmaGEMYufZJ
09ijrqiQoWssXEtmFAXeHrj8KsEdhXBDiyMh+LTAM/S4GCBJSJJJxpMdjHbhAZdosAHBvhW8JGSD
fycGMyKCswMEpe7NtNMmShkhDU7ja0GGbwgEaw+Dxx1lNECgwP45wGjG3wt+jE/ItM1cQJpGZKJK
MJoF31m8Fq/HtXz+FFiLgJs27bK6ne06OiKcp2dGQLReqO4VU1S3mwi+yTg/KSMxniRqusXsuD9q
2/k6rkacujwcsFRSmUkiMO8ICx9XUWPtyappKLi0Z7lAoCZzIvwWOHqZdgif2XTh+L6AR3YozabA
MRbGfUU2QASnhhivMNocvQC5PW/5pSzJquVBuftnu7QInxujXxUwRRwKW05IDGiWr0Jecb7HMPP7
Fm3h3b7wBmp2xkTbfD7BqlAMKJrsK9W250JK8V5N3liBtMV2VUqGKV2uaE5GaoCy3ookbr3OU+of
wS6EfdrI5fehLF6pz/ZrmMNTCr5E9jU/ga7ynO9tsZEAHqvTLgeMnRWcfHZLFpdRRwVMZQKKbAOF
bDZtNugUQhhwpEbcfrdZDXaGINhjeVBNQp3EpV7/HIFgzECRxmyh0Z61Py4YRNKXfOYzFdPE1TG7
UQ0Nuc80grD6al2QOC2fOAS8MLsPowlmHKD/s7RiE4qTHeuMNbNXnVicOksT1GKicdnKF5cVf8rD
HZEgCPglU8xv+CG67RBpVu7/zhkr5krf7AKXJEms3ji1bkw9Eo4zVcWBM0+PhKc+UO89J8PGePZ7
AxUjZPAgmpK6qo9ThFYntxd3cvP+in5aKTJpAJbk5NS+pPtyZfHkqlR8tirjQkI/ELjtLtTtr613
TjmFd3O/3FW3ALQrva9gY1gN/YWoRawsjIFqXtbMjHyw2r2EtG0aPu0sx7WCRsue+KOyOBr5KFgh
STsFobDhTdJ0DyQa5Wlz6hbIGCOCsVdVvgUW9CWo5YTEMG7LodaGSjtIcDXJQSwO+CyqRjTC7HCM
l1d7GJJjjlAaOtm8YqlXTv23Bc6h3Ls5evJa1A2AMA4GObdurjmtk5KnZuEBIU2vD8wZJBPSfCXY
LlkFOVaT+iL+OQ6sWKNljJbUJ7FVHDOQhZWeOid4XrI6488i1brcQyVZ92A4pdVGQ4MCfa1BEJXT
PVbTJ70AKs2m9iAH/dAk9nkhSoavFIz6dGqFibWoafdWf0MC90gYVcJhXM6pwjxS+P11Dv4MvAdE
hIqHNPVXUtUsC5Fl9KbQa07ZOKoUFrM+ShlSct5Z04Fc10C1SWi/7KUZPd/+mmWxYnoK4i31/huz
vd7yWgw19TDcjchi09ZM8/4zDsX7dHJIvNzV8wOHr6E85lsav23Tt5cwgkKR5QFo8xDzxL7WmFM0
NZBh93oOwpDvJnpqdBviJ5ikVcMtWKRWNXYOIvKu36w+O0xfbvKCuY12889Az3OOAayQnk6WmoM+
Wu0U5C0u2Mi9V6h7WVJNj5cSG53fIMC+XyCQqB1N/GfWN8BdmNNqY3qoOtQde4UTpP1sOeFbY3Al
yHbXFtL6kAOhKlsIocmMipsq6a0LULiVY+mmZinUVy+BKp7g+cCltbizn9Tuij7br8cqKEXh3Y56
hVP+w1+Zbm7fOI7TJAH1iNYbYqh0iZi9cFCiqujGRClYSQnd4HslxdST+Z1oPTKYC3MKZDJGzPsh
46/2ndWM/3iejlsde6gLS5QGpKvKoHm9HRTBexgbjmu+J3G9MX09epWltbefCBsd6Ilzwj38Wa6U
xU4Ud+Za31Wv3WGuI2jT/XbFc09aRdw6S+uUWa3ZFKOFDLeXTB1sp8RfBn6OU0RdEma4HwJNNUTO
gkSO87XvGiWq3VTor5TnfBUexw/lVHme5fKZ6QiJZFudJ2AI61OSEh+2a6unvI+N/raYGluR7/9Y
IWDaxYfCdBb7qdDjqbbyp7tnKGYVitivoj6GfXxJ6wwMxp2Dn4pwmGH1uwL+btokJ/xZZntm/l+3
hJVY7G406LQngwlr1PfcbpGHoDoWcy2ZyXXjML5ge2dleXDVbBXc3H93DFQToZ3e25/Ji49BlETv
n9h4HJvDU9mKBP66jXNZG5zL9InZnIRKB/VQiipHq5UxwgP5tNbcDENAzF0N7+1H3PeqKEjnJ5Lk
6UM2+ZUDjq9K75B5ECqX8APDgpNpxhz1ThQANS/ig5KNTw6uAJW66S944f5S0GYfjJIm5MWPxYd5
LIJx2gtDGfpacaLfPOP+78IzMwcFIx3EGqRFZIFZVl9aRD60zox8hSrVdbUZh/UnhtfWwWmSff4p
WAJcOxROE1Wtkrw4TOK4/mJqF8QojfZDM6NCtnVM19yx7YZvjrN3y3vNWx0dMSSUcmk8cdf/0ZOT
TeZfiUDNQqLhDy4ePr/0XLlY4Ed3W/jpgIMAAXCwmQScPBcVGv6wOR5hON1WIm1ZZ7rQBAYy2y1P
jUDPCo9wF1NRhuaOQ4xmbLA0lKduRpCH75F0dxWz/VaGwPaaQTmLeneUpSkAJZO/K7XjbdKi5pcu
n6OoHR5gEJiipvnNAK9Xjd0ZuOAqRml1HtAc4OMo0LQUqnPxEzOQZyUoaO1hbSKfAKOa+u9Yz2a1
qFWGJix7/Ys0efnHF9W8m+nxuJ7iBpyF20+eUYmyrIiA3frSzR86EC9T4qqGYWghOTpA2YK4UUNZ
q6dg91ZWgHzzrjzSqHyc2CQs/PCRg8aQkvsCJiVo7Re8qL1mEJ3Eu2X6lSCc+H5z/DKhBEfaXk0n
njSl/Km5aE8b8rMmCWdxIz1IU4uZdUds2lIXkvAhWNruXGhWkFJqT91Hei+WAG20kqTz9+Gmwhfa
yTuojGrVOaIZx3HznkvE6z8LgVS1L7XGH3jtZ5hktnK9UXOyA82/lvfo7uBtquHw+9Xv+EZuTv2m
WtsGiGKEdXOxe8CNKwtZh2aIOQ8s1SPYF50jI9ukh8/ydeB34hcZZvNoDjFo/wuLi7aRzm71buwB
dNlFWY/yhbrqVe6VJ5VukppP9S2sZG7lQ/GeWrWMpJSmPM57DEHCvwHRoU1Y+xawvFvca2h4vOze
Jxf8GAeRsSV8+WwcotA9chWvyVhiHSLXjiFUa2esvnh9oLqeEB5t4eT4z+O2n+HnTDA7/tkUp82a
5eV0N2PVfmiveuNvrLZEIy/XlyN/JqcAJ7XYgF7FeSISbdEKWT2GK0Ih4M3osObcAmSegNlj7Li5
p3lLdxhjEfDNZRrj7l5zcmHHS2duOvR35Mpq0/brUag7jdM5cwVwpc/jkzQWiPP8am8IPZQwKxNx
cU+Y9K97daRFdYcQxKq4AfvzQ/1Ah2SVFZkBB7KUhZpM9FKDMGSQQV0/PcsCzhbPvToOceGeLTFJ
l7AP2NxuEw43UCDwGAYPHTpUvAlvUVBsCNY0FC0TQGEy8MbEzxcdnyUNCPAU5XeCZlV9Bxds3l/f
6ufPftf31EhNxBsaOJUtUvberCXXVx25UwOu4Lvkp3alfJKFO4BhO2u/I9j2NkfpcfhLXCbVYhHF
+2sRNpe0vmYdfO2/gDQaB8IBqlQtVGox9I4KBufBbQJAXonX4TMafj8iZhj8huqrGQg2iJwoozhZ
BiFJlfaRrQ1sSIHbwS3wUswb8dhZNwTIpNPGN+CKKIUyu1mlqEFGNk1mUTEEKyX0HSxRqaEGTY10
yIpQJQpoPMmchnLhkKN/8hzJ+PJympw6vuQTXB/PtGW938Z2qP5rIZ4BibHEbSLlObCOzGfw8gCk
WW+Pn0xNREu3pcrI4ItyE8whvCi4C7pBqbJsnC3utWlsz1xHkW2kxiSGG+E2/e2ASs9g5q8MIuIG
X89ZfZpGdzQ4QgIcJaiXlmkaRGSTqWYrSui4gA6ftnVaJPf5OjchrB7vJ0gluJw9cYBfJx4WlsWY
fCb/Qs/G5nI531U1/vbeyokWRMK02BX+5G3ydPPkoD0wEDW1JBnLOoYL4KmEl+NGo0k3sZD7+4uT
yxKz4NggoP8ZisAwoda9DGeSRuK24MQAdnI1RvsDByqs0XprD1Uct0uUINqzo0n31pAJzIAAHEIE
HWG+g3Om9dpIZ11BgfYykztoVZQuC9PSgeEILARHoHMrS9pv4bXjWQlJ0Y0JvgjpMWC6LuGKhKW5
rh4seb/pxWk1TrQUdOLNIG24OwvucqVRPE80KoErQTKZqeKzp4mv06UYsGe60xyHpVqgSqlPzSHK
OtN4/hV9WXjlOwIKcEMLLryOAOas6DtgVVbFBjEOdj/YuCdKpShqpSY+tIbhgh/gcDFzYV+B5Nut
URIul8iwCQLfsAMDfpWZS9ij18XJLKe+IRv+cLPZzyG8jryayzeaOddKuJ7o+Hl4uia2f2xTlu8O
OD6YksX4ASkhYUsPusVAQIzNk5OwQtANCEZk1echwysM8OS4N2TgEjxuHnsuhzQjtWMS14V4Hmd7
Ss+KdudXNxWJMfGPQ7I1jZyi7G+m5om49yjtJp8ZcLbwcOvDoeRa3CGKmcNuCDiPyxEf8uxXbowe
BPRCrWpP73njsjDAR6ks93HulNDqDvOFsntviSW3Fyz2V2ySEWXyhMIoGrWhQacAAH9VCQ3+6lcu
cPd/YB+DzKgGbGTbOT0wbfIrE83b5HHHA6vE2ggr1/XBrsdjpHqO/rIzOBeu7qc1uDboa0FQ1k3+
69Pt5MZQm6NbMvfDs6C9cFJsg9nX4bk1To1BPVIUNL9nvyzW6gENX+JIAUaly0iibnMySrd91cu+
oTJ9BerS+zYC6eGvxIDfDCLSc780fWAndPw5jsN6mzCH1H+boAuQTGbqb9nPS7DFi2YzFJIKNT/B
8WxFFj52QT7/ZLy0rxlVn2oQLHGa8xHpXULzVxyuSwrqeBD9McArpOLh/5hk3OTImRkgGtb2uVYk
bF6/StyEGc7pDrIjti8o6Js0M9wFZz4Nlm6NeXN03PxO4T3BBBccDhBYd8oFrOblJh0bQqub9YSQ
FVCLHMQBILjQKtpo9kgMv6DLskFNA4tUHjZviV4VelXZOPfBaF30P0ZFQtJVlFZvDW4eBN1bi1eM
KnjWnJA8nVZRnldttWnmH3cV/0mHXjwfBPvBxvij8nDN8CTqiOgQ+/xaUEVSgJbQX9M+iSXCpVdt
AMDIo3iYLkmAArDhs4Tt4yKA4PgVDnhxM6ctwvUI522lTSTJpOfAwWjxMBXm4xgqmAKtCxWXf2im
T7EWqBpegr2ILtPniYB+sV7b4syh46L3f4h5Qjy+qLesVlZoKl2tEKVPVWXxrfCToAYpGN6pLTMh
OnaIJycIJayBwTCDCcl/1KN6xNj4slLO0bpKWPrvsWrhR2R8eqwX60XuqL2R/B8WSZJ2HxyZayWL
EEebtbwA7jLZTN9rNIfH4kncQRZpNeeFIph2r+Aih5B3U7eKnqjUnsxnMkrbOtLrtWCHte2txh5J
dj/t5iEbLyxsqlvU0hu/KkU34dAfuFrIitItnWAxrtoslXLXOqh5yieQZcEk33GpLwgQfkASoCOw
oWAyT8lFqKS0vFRp4U7skq/eYLdjxNuS6jbQjaf3gnHONRzgEOTJylSULv27D2/Jyc2cTaHdAx0w
3NDVS+BkrJA7sCJtCZniE+aBwyCwwOm+r5w2vV6SYq3yVIvGRlLR2Pa+0hzuG00aR0YilHsfwh5v
nl5fWlBtQ4VmlKZShnT5ekYvwXWJ1FgcAcQVGg/9sjv8VHLX8a+YlklAryCbB9u3+nrDcNtz373W
zXnMl2Ik4PYMqbNrOFnlyn/BZk9AdaklcblIHsGyze6oyK1nvN9Z6VhaHAkyvkA6J3oIoX4jGHGj
pEdGOrvTx86qkn1zetSjCgNkZru7V+/uErurBlkvCZBDq+LhcDzsFWALvwSoJDXKtns72q8UIwZY
uWGs184SD8FafjZFC3khjR3EfZgjXnZYKzMJcfZeLNrPHvMhnHsYQcj9YzMKXz3wc0EVCAaGllN8
eocHiiDcLJ6cENwpTvGNjZxu3KtJhOb2pwr9/Ixymr8hD2OPNnBjp6dunwnsq6/gCYmILVPmZC7b
NCH6BXCp50HqBPwuN8jbCqNm/CkEtNAWF+udR3KxCOvJzHjJ8M0CIFHzm0enaj42RIK2UtmeGqCC
EhJyIBDSnBN+F4EbBnuW53hpflXtu/XvtSkSfgyMvc9ZCfpSRadlEf+3gkLhVJwoMBAWEJA5w9pg
buBKPQqO9jkRbTTFB4fa4KSMuv6eq7/YQYe0pD7lQwh/rqx92nrQBo8RsAdqshbmAmZx+YmLvWFN
INZFg1zdNmvvxvd9btsOCFvx7AnRPtihFnFnsXSQWGiGPZ9nkPkT9pvwnB8pFQa0b/47T86DofuH
xfCm+ziEmjgBCWZZri3MsazjNSsm4NWkjhCGUMTta1rj1WwpWMsFD30nBZ4Z7rq8uQTSvqOtM+EF
oSdqyw6FRBOevN+PfoF4/OnZVGPv3GFEt6W3OQJMKr5DsNAC5R6H4Ya/vOsLNU3F/+H227OEGVf9
S/ROPEaFi+HK4aCrOhZlrNTX5BcDrYrw8bZhKb8HIRCZRaFFsqBbbDJfUAa1tCRAAfuPJe5I4Ryc
vxuHwNrIGgaLjY5YYuY05NwcV0TwHoOFNfawmmjobb/eDJXV+T/mXTTFfuWVh6GNrkBTVfnCfcdW
x1vdq/5Ay3Lyz6RTcNzKdGco6qgWiD4z7XsyGPdhrrnncZsbR9yxnNsoQ0PUPJ/Zn+pnBJ0+unyZ
54hmeUhqIxNPjDwTVTc3dMaRB3FxwxX/WYWL9IH3YN9Jv4j0WWneK2eRCNRcLMGP4SEC+UpvXRJt
Bw54TClX8S4sEinMAKwMnQPLYaFLK2Nii6NTW5aCBVaF2LijVf2+nm33DTj8uI6eE4Sejey3Rhkd
sta9AFhIC9eZA0p+Q0DB2flar2HNRQYLvhfCSIGahGczA0HRv0ChIHeVBZZHQWyDy/NSK6nam9T7
+cfEgTn4j5ee+majq5j1k2R6dUnWQ82ChCYNo6o2EF+K0/wKT+fX8aEzY93UVTU5GxSnK/UJ4gPw
fK2iqSTqETStHkoii6vVkKe44RsyUuLAUW68UNBxPOaXxYSmw/3LXhKoemyD3133CN4ScenZgvUg
gWXOZrkm/tcYqq5lmGI2IvMtnR6Zen4NQQbbl+85UBUzqbvtDs7y9iokZne+lIDKzRQA5qIQ2CcL
WImBd7orh/K1Cfp5aD/mezlY8A6XKYHZUC6ngC0515wQkKQ5rdmGYwyyJVCBx25Iaiuyh96wpM2T
/OYI9QWbdzIJMeENIhE9lUJrZoQlW56w0X7ofXQixxVb66WoeY7//z4uBhkiekpUV5wu7QOYraqT
x+G/VGKqh8njTrzMkALuehiEezDXqAgqavEcLkcKJhWiTL39hGwmu+0MgnU+nTJoXW6HBuNyBaiZ
cMzwRSEf1X0RV7uE3JvlaUn2DmDcBwGhMgGQhn2Za0EjxzF4u3853LsjxPgdr4pNZ/Rn7/Ic0nKs
d2TrceIlQ+HSi5wA9jJ42SY1Ta3J7uUF0if0zjj2l9H/du8znKLev6xR09+ZwLqCaMQI50ZqC+Q9
ojFYNYjdi4FYUGPecG5P5GxwTECJZfYRoZNJP5qGS+03hbD4akxCvaT644qv40q97Z5bR8xpOwR6
FHC22iDANGtX/fY9sUiQHqQQyz2fq6VHM/5pAdpRPcX0dwEuKTc6l6NZPvjTxVDYa98ZxdXkP0A9
D+bS+fBt1o5ptBRkVT1qGJskw+EGCwOwXg6nY4e7h145faJZAc1MPWburqE2MuRssDwFvjPyd/HM
qWAuxIzzRkabEz1QOsXrLVP/kZcaGuhZ1vUjvFK72ac2F6ZfvtO5ECZdkGLcepZEwGjTdcmRD3Io
JqH3/2ZEOoxYVJ7T6TknjgEGZMAj8Nctw1QFdFTtcLz0BfLZlguFTmt6fHe5Wp5pEwwIMoC7DgpK
q+Dp4++/gtKeq87cJB+f5Lzvmu/Wc05vsYOc7OaaGUYErNswUIIvg2kq2EOp8VaBHn2fmqR6MT6T
tU675rXPMJJUPnnd8CYZ7F6bdaR58HeZAfVzkm/vBsEmFF7LU8v4q2xqJUkxpQBvt5s6XUIhlN37
RVKCWmAeY5ZiZXdwHZYH5TiOp19vVEjNn2VUoc7e0Xyqm4S6Xa0eb+ALI/GNPQIrmiNCWuqQXGji
r/9uCV/ZTEoCn+CPrb1SygxQBfwMF+DVNzNTz9p+CJKKYrcYW/rNHgSasrWGU7RxCVZqJgeZzQRK
ktLDXPuLXBJzyrrcqntcNdy+etlrlH9FrmTUScVeQX9cJK2wXDeDJU+9+rdAqnq+0dFEpag0LWRB
nZvunsgSVUSHVHPSWrB4A/uA3nvjW8AVd9kO82P56cPlWuvAjnGoE1J4A0gNHHngMCLzdRqP3p9Y
zC4KdrXdTBIiiKBNXCrGVwnfvSf2wGgKVnPmYW8zwFduYdOYgotioSBJyNxSUieY6d6pV3goNry/
uI5N8YvxdZJnlPqqRTTmwjNIzXLsULxX5iQZ7yCXIsgvJ7+McApUvAruM72+3F8cAfV8Uavk2T42
xY4/t8ue25tIiaySLjfgd5jqE92TyWxuBr/1qBVgtdnm0/3ZptlUjFs+dGXi4hSMp27pHuhHfiNL
f1WrFzxhbjkPlTfiLMTes3/G+9zNTZ1WcAtwmHt8FYg54F2w3cCZKnqM/5JKxkKyts2vNsS2C8vf
fE94T04hr2qc6WZ5ed3fn/cN8ilRaMr4XKu4QwVHPoBv1ACeuxdEryYjtCLWAkc0OG/eRvAi395k
I8ZJ2+KrmRTq5YED+d98V6wpGXBvlEnm1unbKIqGuLquang9iVMkpWsUrxBMdWJttGg5fNVwluID
asrIGaY8ZlypafiHe8LKFRVuA2DSFfMsICh8h7ZWZ1rqvwz/a43e8l5e3JOvLfhFF674S4tpY9vZ
s8knckz05JThEaZy9ijGyXhLfek1AebXncvw6Hdmzln/MfPaAKImEPeL96VObTJkVBe3BBiDZpZs
xVi3Piq3Iq0gu4a/0e4js5PNLSBR+wIT6pnsVmLx6vOQ0R8DQYL1wWX8Nyxjb47lm8ecZo55M3gv
yG+0NsL/f7jhH+1PelmY1cphqtpBU56Nbeai3SXiQSIPHD6ZNRgx8XKVGZvwQ71sLfvSh8Bn3UO3
9P8KLLqTBCL9oSe2OdrmNK5+pnyuCpJ3zoV6wzDXK5flWnTaK1JGn5hPbUFnwEkgSAuV/A2Ny0vi
RZKVqlLD1dI9UektbN3XaaSrO+mK3K04a9P7/QaWuVdxbJsD0NlbgHbmbjbriuS6pTYqo8iXvDoi
D8ydtawMySfBST8gnzB2RaBAO51xE7+ikq54GgBOxnGDgSkiKmd/Ivz/DU71Yz5ucPZVUPSTPklU
gg6UlPNXhMWaIBA2fhJyUTEUZhYAAr9VA2x2McTjt14JpY02gElbDLJeBJT9xWoEmgACpHk8cXaC
SrV51I3c0ripMKrAhBLjwlgY4DU3dr5jjualm1u0NCloMimVmmditFhgKvr2zGSF2gxB2B3YOWLn
RFSdVJYKyODSG31lb/X1xkoN9YjbQAV+7rLoOHDSKxi15st4hF3fHu9byMtqTXOxDIlSLSQCxSDm
xJwgqtyw04E/5KYb+xIvk6iDxpJvUNhnYfJNYbbU36iuirZjw33nDwc2WgQwFIKN7cjFo4ruOATx
8d2ipSMGoE5o2EKZjd5kMiC6Wv5yrPSiJnNZuxlqFVBBZT+X7NLDlX9/Gazyo5LUdAggxtUjDaHA
QCB2bJ55mfv5U5cyRF+o4S+qlnmLjZ65j20e0AE5eWTBGkEjxdVOX66ytBsvQMv+lHhYHjlMy8/t
nkEKa7Ynq7a2UDD7RwMs7d3c2IyycxhuGkrmDbRa9gWXzxahhpy/0j9NFpzEtT5No+5j/1hItqUy
faXTwEul9b3jWhb/cmiGPK/blDfQWWKOxxLowCkYBgQ0gWZFDRuz26BxriSZFGe2pGREsBKz25kx
1ML03hT9aMzhLak4zffsNUMZ56ZODoYVYBVaY/nAmWn40bzFyv/J6aRRNZeIPDmtRcpW3NPvfTCU
17JoBI3lvMX5UamIEfnwMpp1VWUwoAEEGkgKqt01bTG2rrT7nt+vQmNLwHrt3wbqFh6Cw9p0NiFp
KsUWIhPUZXp1GjEvhZQeSLA6crQYCX9M1Ut1yMiZ0lCl6CLiuYzbf2/slqNqaXyjY+BYfp+FINIh
a6dbFb2MsvtCl5vYTgcR7OIqOD8zmWuRZF5s5bccZfnIu83H1Bel9Yj+wilyyX2cyt6KA5a9DvX3
teVfZiYsdexAuy+8YMmw+msapl8poJOLL+NaZN/1yhf47nXS15fR1arQgCP45MXHCDH5t/XNGP1R
SJsTKIrFq3Xw3gZ0PSiMy3Z2VgiIWmB/sip6ZOAn256EIm6XP59h1mI4YiKWnrp4rgICNKB5iPhR
r7UJNvoxyQz6J/5bYQIy3K2dteOME4fwdleoiHHtNQJXkYzes8IQvH6U9M+bfHyXbSWlkLGBJlDc
uBikHbr6XtzSpmhelXD8iVvfXfpKTT1EbRyTRXmQODMU745+eOj7n1O40ruvwkn2WczwBF+Uv/1b
tjDPOiQnvMYY7QarOOwkHewyit6FMpP5FcH2glA4flrW0nyHTaFQFb6kjiJqJXyDog7YEJA2Ecz3
5uWhUGGycxmDtTZVJ5c1Be87taGSjq1973mjb2kd3O81sU3JBR2x1rN0N9j/EXiCaumJVt7Bev1p
Qf1IEYH9hOu73+s5EVEKRcYdM2a/TjDiagR+v6IV0NACdrfdWEsPL7iiV3lrmA8zggbuAKcDdzQo
x3p8CWlJCHzaUh/6bY5lionl29ud76NasZ47waFuYWDIsq2KuMalK6AvORfgg5jv5+w/oOW8M9gK
Ag6AF/m0boP1nNvLQuzFPC+675Jg5MOgfs0YOTNJ6ZeqRtMx4c7dOomh4+YQ5U7pImGRV/2h+fcn
EzvhjzjSfeusxmuiMRQ+BENfPkTa/z20QM6ZJZjRDOcPN13MLEiO+hABLLwXaF5YqpNoWFvs/ymq
YAX4mYnmPJA5WoodE8gk+dgoBnzRhXDquGavY7kfcg8jyMws+H08xfAr1qX68sQS8BNNHWXvIdOW
bz5JzCc7RovWNOjBzQwUKHXOA7CCVxvAMNRia+/CBnCgpQSdnOqdk2SJs6Qj11UIYEYDpSR3QWwu
6cgm9JT8P0L8/1zZvKPSthDnxGwVg0kqb+eChlS9DdJ4rjLUGX8JlAmt+iWQaGzZj3zEYjtcIFr0
3CHYGladqXgJPHPtHLYRWCqxVsyiloAr9achptaAVvX97khNjLRNTFPdBumKXKiGY6vnVAKEG3Ya
16VERq4wjZzpLT0Xdh96C1fzq7Z7Ag1GFHhQ5DOa1iBEJfiU7+F3DTJyLSqajOylKFFGJT2Xphd3
n0UZRyZLJpRUUECFbNyFgAWOfR98K7PEmClTtBHu54BIjmlYs+J4iIWIP2Ep/mCfL4+L7TIzEKis
HPoadNnDkjl4aK4aM3Tx+BqeA4bmk2CP0byJ7hyct8OQ7/Xjvi5hTTtTRMztcDgRxgQBM90nsSJA
sgsY3CNBgV7jMT8lp5qLXAwAamVAM7In0omqgZPosjFxoGwPzOD4/CLsoeSIuvQF2LZvDLHQ7kem
oS2BW54J2y7cs1TqdGkJbIZZt70of8vktm89tQ/y1fofgzMxNVKl7zRmvqCPSwUJdM844+dSe/cB
IUwXqRsi1CQqJTA5QkPYj5QQUssaTkM6l/iNmBykOYa23XaOZsvn0K1jns6tmOIPG2JmjEddWiSm
/H1I8rSQjB4M1HAziPkFdzBNXDrJwWdKsYiEbgZFXB9GBk8cxiCfTZnY9ngjgVPnAVmzWgUa9a+l
wsUl57T/8GJ7Qj0IKelihA4zxX6Ef9wpO9Go4yiVnuHihdRxW99qQueMJgFHKqI8pboSNEeyrhHD
ofLudlTd0gxIUw28oFTEumlKcdskqHJ9ogusCwybe5vrE4SXOoLi050qXepHImT316o8l1D6+ptd
qM43vKL/epjKX1IixwaN7XE4hA50WpVdw/JDx3K9G//d4CiiZt+XUQbll/7N4mPDGVqwpVxlyaTA
1XLxgkHVJKaCODj4QbezDQpKma/VcUvfKsreINGjBuvA0qWWFYMHRPpJEDzfM/lNyDhfPd8mbF9z
B6yp5lbR9Fmf3mJQluquIif6pZmQHxVO7ZwFXVJLbQr3HbfCSHNg8+3BxiNkxKlWTU1eqBCCdy0t
xWZ2FmpIx4s+17tXA1mbPWU4Dco8YvK4zegANXah4fvrdsxb8hLgYqzh94/kllGt8W2ZGZaCzcRk
56PRSo/JMm5eQaeCNfaYMhdzckpMfC2Lu+G+9lx8vhM1MTNLO8/zpS2fH0iZeMI+9DmjevvfdjgY
6PWHSCgnMUauZWA4MKRBruK5Lje2BlsySqSYEkT0f/463rgEPQ8Aj3gYHQVs24uzS0sFgYeq4EbV
LeOdeLJA6kxU+HvzCF3rgG0m7sdKD9ylPC1Tkd1jYC6sOpIUVg0+AlNOXMy5/+C5z8tv7dW7c2oz
QKwf8Xb3HGprpYYyy9zgG01Qj4QAjJ3je28X4Kh7b9d1BogxQQtQYZb5AMTs6h4c+BJN5bBFlCF2
SY72P2b5Y39mDDd6iwkvqKQBupD84nuFIzfHu5deBX6PyEZNrms4A1xTSSwMzPOOWSuE5FV8vzbH
v1pfC0ymWRljIDWb2n8efyPh4iv6MenW95K8AwdMl5wMmj1dKIGZMqSr3etA9M2w+CSgoZ6VBjHj
j60izWmmCmzVhTwP697s4TlWLEf3qr4+VK0B1sr6TzsvMm33zIr/FfIEg8R8wpKmRnvOTHvkBZNS
YrgKfK8ItjaoPxZtryW2U142s4MvFrPdlTC9u6egYP0NKT8McOGiMtCvRs2jCEYba0dJHwNJasc2
HsT5kmEFScZ5RGpCAuzpqUXhvOWLIwobc7XfuIN/NzVFYNZ6Y2OwL4AWNmpqBRV0r53S16Ddi6sr
KSmwVwSg+sQVJFKZWn9mTID1Eb4mEJ7Ypbff+b1pAyliMVjedF9oIZzk7PVa0lT87FCXdWHT+7WA
phcM76o2ZwKkFqv/W6qbj1JwyK7i5PEeljiiji3djeZKm0TWOPJpephEjrmWhodTSB/YA/g8wzDL
MYEhE6weAsRE6rZJPMCXtSl0Nzge9sW825y03jp6xqWTuiYwJIp3QE0fPulb21kIkpTfubw2rUkO
KfFOR+C5o7XnlGx/yu9/bxrw+aGI5H9HUWPq1tyLHMwrbyQyT06/+IEyyMYc7GvyRUa3LD74B6WE
vpFZ2x8Xh/4dyv9VmNe77z/zemHq7bEcK/uUlX46wcxDYLMoYmuo0QqENhIfKNRWblPvdc7d/TaN
c0490R3N0vlPTZPWTjk1ZwmxzfnIuHFfNzhtC/3jvNejdyEFLhO3b0yw1zsKZSeztGCNI3XnJwQH
MPv4Ff2+uQQ976s3DpY+fE5yCewZ4t4ua8NTzZRoayqaARfv6bJw92qMvfqP0I8tpSaXTIdDmb3o
aQ4C3jRrV2teIfuyurxnR6j803gQLCQny9AFfiiMkqv4Cjo7b4d4dpZ7DPzeWFSiBIimC48DJl7c
FB+V/fiwpiZhJaTdgDPgTqVvrtdWVMX+NbJZyTrm7nB5RhbdODQ22FqqKH+Pogut+a1lQ7Yjc0e8
zSjwcT7sogyPYm4eX4p2PRnTKSgvLnX45VWgaun8zkt9A2FCmifZboVtQk5WpxviKXFrWeJBsvT0
pEldyqp9J1ZN0PEtALZRdcH9DcIXIKd7fylLNlj9P7Oi1RiKE431LQLUvZtJXmJ1cnBU9gOyYvBZ
1urJh7zSpzB/Yqt9EM2gEd1NBYdM4nKAK1VR1uBYQjCc9tkMKWQ6zUMbzFiRnxd97QzwQ0I+h8to
PYppQ4LuVnD1beHzI6LZ73lgTNGQp0/dSLBOJnGKBLdDV4TlLvLjtLkw7nIxTO+li6KAUKdGUnKc
zYHkeY4WRWrHIdlo3pAP02wIO9hR3A1NtpO6CIgdHC9+js6852uCBbyA3LRCeKsd/nJT+GNBDevK
SOhecvsMEVEVVIufMu1e7+gukNJtfd2gmmzT+z8mbPE3lihU8HhyOy7xvc0VpTSNcJNpsFm++Dzt
DlY5we+uctAW9lfmla3XhJVVsr65fdy9ZUZCPoRkPNhAlG4UrksPEOPXar5Mu4i2Komjnhlx5MqD
sP3cV5jk95D4JKpCZXhH/JA82v6Hj8XVArLwqq9ua/skcrgLZ56F4c66eOSTZ83skqrTGDsi0f+l
pOsFisJmw7kbIeMGhhZJcupLZ9AstvOrrxr/Bl3IAf6KzNezVnXFZ06MBfa/8MGeyCU1tHHunDvW
ReIqeT3zDPU3W/VwIjHN04jhYbOZeBRGFkQq0aUnq+4RbTcaic6rK/yF2W+edR1e+QWiJ61nexOL
1STmU3kQEfRMS9rarpudN97iNxCga3hah2hB67vlgoOTQ6RNWW9eWEIRGyO+Jv5gBXO9vihch+uZ
9/ieVvhBnUvQEIbH7jPUfhYTpU7vvno4QPoXp2BBRcBxudaT4607xyX2TkJn/deuZ2sVeZB4BVix
vkEL4TV+dln65vCtMKmkPhK9XmVV4MNR3ZC++L2o+lmKvyrUalys735JwENma/rHRq3x1xuZX43R
fmNn5N1UMBKEGeXAvMPCEeJHbg8wYWmZy5KY7LCM7Eu9QW8TtKC1ojQfvLvFI+sQvQezul2GKH7M
NThjJVFt3TCuwrdimFjfRJHjyxNkmwF/BswubdGAvhHvpQtBdwlrJTDlK8Z8Bwep6T8Hz7Xzmswd
oYdkAdjCA6043wdoIs3xHTuSrtb85RUXZFXlxIAYIlb5xUXfMnjIWRovh1405F1wCg293B+fh2sJ
JN6P964L3YDTBzoHGXvb7zXkb3M11idI8EBo84dUNYx4G3k6SX7cyodDrccC0fkKhYFlH9mkKHBV
3sq057L//mm7GUGQyRfXIFbBamR7K4g4qb0whdllFEtVrrEg6aSzH5Ki+cgDAsO7SzviML4R/Tej
+odkUq/U9/MsTTi90+MvzsfEzBJXFFdzSfdtK3ArhSeFXiVR3az9k9CtPeMvbOCrgkInTAlXSg9S
urWqKAd/IMePUYsihaWjhvNutrBJH9pLT9F1JrHk1jEncixjOayuEo/cMwMSaxAhNTbf5+IRaIps
+Rltrrm+M1xF7/Fi45MnoEexT9crfxce8bLl+0OMqo1rWonuInsul2G2HwdCI0xXMp9gaiOLSpOX
c1MOHvmciK/OTDzDngacLpPbC6JS5iMhhYTTe68TjfxvCjM4/TBXNxT6KoTHsTGpKHAmkhXv2paK
IkIQU0m9vDD6WlgSZ03PgdS0U9yk2QJ8pskk4h0+WnJIEGUfdHWSgRyezNrG3IqY27u9WQm6rYWC
1Y/D0iwL/lhFOfWE2+Z8liDWcxem3tJKn70bqm8R2PMXsa9mLUw2+uEMBJr++zWpUABcQ+bGThAZ
WpdgV/JrDhOAF2rj5oF2hAPVTnI7hwbs60SftXXtRRGBX00IinluANe2lKShpKu5YlCpCY8S9+TB
2xMTbr48EhDUHFKBpXRKlzC7G+0u5ZYSvp4mKasPN3aYKFSEwJriGGdiwpwstLKQfRaUjt93NMbp
NuRFhUvViU6f8If0nSLHUZwVr1QQVnuRgfiIlV9ZaPzRXsbRapVQVF/Sqx9sUptMAlt1WvtKNyF1
hmnA1hoaO62oLGuPs4BewtCQITAgVadjSr9CnrZxB3tqMf8xX8Vce8COFLfyQHlJbCEPJEHMEUaO
cf78/dxPK9r4oGklI1GCdMJOWNxxXLrGyECeNndUEeq2n+1CyMM14JhCNc+ZL8xSKfw95d2SpTr/
eQsW1LdrX3SpNXG0KR/4ltunbFkbMYvDYsotNEc73CvR9sBYVDknb9xDPVI1sl9DeyGQCy11sWXK
FJTI7s2ORZUp6uBYI2NZwEx2A4FFgV5pcQaUrds/9fe9LIBLNUxvoLZD2oYvfLINkR+YylusKhj9
2HFU+iauTDq013FMwVwLvXVRcmn4cBj1b6VtmijPCY5Bfsm4c9TrrmIMWs6XqHXednxNaiPa8J+8
xyn3lGI16Zkx552awISDzxsK9wLVrlkvUYEDXIDyzV08qY6mxZyE0f0nsdZ+MRaBOWp+SSZuHsU3
4hbOSgQ51BSNsitpBAW6mCKt28gor3vOLrWJugHDWlzufyGXsfPSHFBaWKSPbrWKZADT8egltoNC
3DVoT01joAYCXeaPwQp97PliqZRYD9+85+chn4LLg/WhdQ8YVVecAae9LQyJjheG51KzIjG5d6N2
7jovtKxV+9KTjW+iFSRNH5o5nxlowWnVT48x+jemLNj+9u60iFqOTprfkXtrxhkKbctm7sc+q+Zh
NR6zWPnv2SeKVwuhBtzlMzzKCJ7kNDuYwCtU2CkGlsV0p7zVTaOUtC+jkk28mHPrnYJx9bsbePFN
c03B2sghmufvRvyh2aUHO7tzqVcULwlQ6miq2gdqMsiRxl+A3oAaKg/xlLQ85d62Gfty4EtdDbpY
Q2/FQ2JZh61SZm7YNBE0rbwWkdEhrpPo3/CxO+GnLHzxlzS3Kr1Z6xqdUNNXRbmSWgefWIjmLGo8
5KGpPbazjtkB/m5H/bUaLVF61OGLYfRcqxdRROpkn4HJ2+98/bG6FLY9qXCIBGii3cgbF4Pq6Ti3
LK8JsqQ98dJnSfBzZ1M8AaDyHo0MoWYD45OdBHK+Vbh11QtetK68mPY+KJIHNugtmVxqiMBINXbu
a0scfOhrdwA40RzRF4rCGGzMNRic4riQ+0ULoDB+71TCKG7KhEk1sVM8lFtWH9buRxpienlpJ7+N
+t9/CLlGIT+aIIVWrbd7t7cwz9LcmV4M4qzLnbtJeCwIfPzQ4lIRoeju3YZQPXAT5E/dQOnH5npr
fmPgzOZRTL2Oi4d1G3+2jn+4hXkahYe8KYRxTcoNbPSuyZAVOLUnBFqXYysXtZ2oBg/fUqaW9I+6
SgcINZUhqSHTsq13CaDre0Wmfc7k34vZ17pf1R5Op3mId8GXXOgjaf1plA6bMSD3+mQJ81pCs3zl
AQauV723xfi2GYU/du9ITt/LMYSe3Vh3lVe6fFdoRzvWPs0T/T/XEPMEPM/Yx8poyxIy3OdEpAS5
/+NE0GUM4CKgQvt/cFZnBOwKrP1OaUlAz4zrSnbkgTG3ACzhENnq8SLDSBBfS4F2SMS7mb3q/q5X
f7vbcOOhGVqUpTSvVuqDx3n9eCSBRQgoE68uiZ6ONzsUIVw2s57KE94wqI/SQK3enEhD9QJ1B6IJ
TAn1THpm+m55Ufug5pQn0sE+BVxz59F3JEqaC8rJbvmow1w320J6dJOXS81UjyR+RvR4X8OqhdAg
BTdnYmKOSIJLhW5+r3JzipqWwSGXeiPEHoEorvb06ukqDXaZmi/M9Poqh/ydIGr44dIST8mrNExp
/sVD62Y9h2QTUTJGj+1wy+Qjwqj1p2DXps407yZTcsY8a/WShl4qLl3ipDN52/DHxkBZfo+GJzzw
UiNw12mKapJIu3RIoVy344tLpJT3dE3wB7N61YiJ50q2uCC2Wi8ZQaWnq4F6jqXe9OFsRekpQYpz
gSZHoZdabHZZ/2vnSrNg//ql9P9/SGJgdZQfRqD3ZMRg6T5XciKpYOpReoPrqRHEjtthLZSj0aMQ
YwwpfJKA7UJ+OaGTETCA3k4bkiC+2pUcAcEqNNimksWEJyxxNf1BHW+4QsJDlXyTOvhiqVWCOtQ3
mV4vSQ2UIT0eRWyVvq2+hXDqFNrhjlGpl3PizplDwDf7a91VYvU2f+zmYZ7gP2CRHoPvCU51+MB0
QugN/QyrhANSFrTqgzeP6rMbJ3IjgFryBM8Re90v81B5vjWXC8RJ6aheJ3H9Di7/7fl7PtOqxE6B
5clNoVpvLjqV7raLfa3Q16QZWiwlqONCjKiRqi8AeAeNpPBqZd8QLyh+QMgCVj4AVouB4til+FmV
6WCQEurGGf2SUoXlflufDc4GHBbSe7QWuyLnTPmEd3QuAHPIn9jpXybyUuq/nORYHV4fVcWr+v3K
baOlU+ConlDvIloaoJguNA7xpl44QOC1EwQt1moPmqnkBt2apb6yhUdOtptge8ncgE6qJj8Y/ENT
2OL8TFOrRrFjt9jJ76yzqWxHjrSZGFo8hUZRYb/8zGfQoEeAd5UbhicHyvJ+23RMKWL/V4nc1lRV
4dXkxNVHTGMVQ9CZ69nc1Dbzs9TwepdngcXPXIt6Lm61c7vPUOKL1oxCa6BfFmvAdhYWam+qPer7
Nu06aksr6yj+IpNvWRhhcKaSXmFQT9RRFD67tewmrrQYPWbRW7Ya1KoWkE2/hLoFqlvVgBmQ1DXS
aCm7aH7MkF8vmtcRbVxGIPnN/NEN21LQRvoFFWs48u/ckJcomrscJ/bjHxL0htbdzKRS8mB+mLen
JZwfKSSIsiCSQH0ZIXwGGbZrPsoXLzbNCNpU5eObtwLlN+N1JrjIT3yOpaGuhZfVfQBl6rvyFoet
KIoxAuWyAuJCQB9bOqRztqgr/ZGYvLvMhUwtNomukLLsSZnAFwvWchXEOXkhzFkYah5bLzhkO3hU
nKqWHZ5GD2769heeLg9D/faNnp46X4WzkUzsk/gp3rxfRO9ZLt0MnCJUOlzhXLlpHpvmy9Lc5iRG
WJ5ksoFK3Zw4evaRaxTltB+F8b2NsoxBkvgBgsn6i5mKScC9BhsiAXBKWZKlu4feQL9C3Q5GnDbC
9DwkHZuzEKXRlOq5v0ZP4ZSO4Ysn9x0/Y9pEiSOVWzwT6ETpVQ4INzZE+OZsQlX+ApcE7YILB7c9
cS+9C5YuX0ruPL88y0uNgO21juRKLHhAlRZST42J/jqqZPJ4wXPNum8WyJlwlhyVnWlVP+YtlExm
aTosTnPQg0+YQ+mbADCgC5k5KtYcR9WeDFClkpa6H0DnABVyuD9IBjfzg+fZh7R2fDPgJlSeGFG3
464krQJpmS/H1ZkN9Zf6r1YZK00r32LEK8wfH6hvsKsr1hYGfQUmrpUcTmc1dg+mXKuQZc0QAU4j
+6BiKe5bxfb7PPuvK86vHzoMAJnWgGJ9n8wTK4jAvAWlhuSOViYooWOy6hz8huR4Wfex45xzsVLr
A+dpJis45fRBU0Ll9/EoNVGu8mZNBr9UiuJNChy2AhsETG3lcpmiGh9kbQDw3dI9A4Hn8Woz9VB2
Mro2YUxZwM9PS/2WvfW2rLumAH6UJxbYo6uR2CrQLsuAZxeHn6OIYHaHXDMIeV39I4XYydtMw/UZ
8VHEZZ6hxcv/Pns9jLyCZYJ7frHjmhJl/qZeotQWH3iraGouoUEzDPcdYnW7wok1n8HudwMnu04v
6dyt4n9xgP4r/AXrq+HRJXYSMcs1VndFnNPu4AeMvXifXXhv0n1meNJCWvqvNKVGl6mvTQXE36Wp
YFf+pbBLAbV1L/4v1y6GukOM/Dt9kwec3BIRTYFy3pehP+Y2Cqr5eoFg5FdFZ92vZ0RPnZLVmvOo
DNdG7rgnPVp/OuPLW1+duYZ38BZG2otBVBO4/01a3Uz+//c/1hZZV03Y8A4Oe7Q9hShHINDYGSWg
TEyLO/MZwWuFEIQ2ep4t41NiEDOkd/iRDi3fXZVdnM9fjuatmX98QFySSZCuK56VtXZ+AlzRSUb5
BkvZoF3VrijTnbyxL7zsV6JTVCXZvw6oot5plxIg0j/QGz8fFnN6pawdebAMNL89YS38kjkg3et2
P70gJDy8q9kxREcQnsv5xPLYfCdICTZ2yplWbrnbuD05dQBiyAA1Ra7h9tYE2LXZG7AxKdyNOAyV
t7rsjyAltH1nELNAVO0RrHrE4Yzz4KuNF0kYESdqJQHhCbES5k+9J/gmdLQtRt8GjeGJ4Y0jMvQ0
9iusm51fpG62WEAMavEUqILvvV6jcKDrA+XPMAZQNYtLVnmmH/UgPcDQ+xym8Z7r4jkg+OwpAYQN
3gE1L+kMoluNoirjcf3P48sWHLOua26RxjaoZlUUwTD1mFDceeW+TMuh2dxgDb4ReIV+J1mCPO6O
jgWLr1Nh0nAYTWQhVmCfEnxiWQdbNqtpWcohKewP570NerBWktwR3lpNq9E4z7PzqShElbTz5Bpl
5OhmgqI/5UymO15Gc5e3DK4EZcwVM0yWnl3qRMQptcYrqyqg+wZlfGgNBjz2h940IWjVIPMJN7XJ
wup81khOf/rzNktVDqkEhRooIlfAuSTL1GsDLQt9BXl4p9WjSlXJx2/JH8FyFVd65EDZRTjaodOO
0tABVaZgEETnFYDL4On8oRoTii/PW7IAANAMJ/bvuYXHPBTQ+AQXfibk9U53WtSFHkcbCVZApihj
oShVC88DtEz71bIcYH0Om713vG6aROhH1rHkQZftCutQxhEVhggaA5mrIg4tkF61GcPMevmHvcEU
aaQOxYM3OouvIBLq4LrMO9jyif/+2x2H8nJ7HqNyC7tHWM21ewDI1kaI4BuSAI/s6EIxl+YpZoW1
lbHYJAPP+GjaRoasWMbJFw3RAY5FKVZ6lJvAcfLv2z1vdAKapLzK0ZynMmlMc8Q0QAmTu5lPNjj9
ae1fBgYFqhY7LVTX7cR79MrddJQBfNgVn5kDbYhRTFtC1yWbtoeiGQVgcL+USiJnDewU/d8G7S7Z
Jog0H486PtWM0rjRDdr19+Kr5FT7oWitJYWnnQid4fSPveRPOSDqzWLEe6RM+PBEl6p8TvU7DZ7q
Lz51xUx1ZKIOmyUmak4Oe8dL5cSu8zInPLnFHt2rEVnpG6Od/Py5I5z0rAckUQWJrAx0YOZKLqhH
dIhzDTKW3nlNqQNBp1QXtl45cb9FEOUMJxZcvr9PC+MW3yoa0FjEbHyRnsRLJ84jWQP8MTayzRUf
93uRCrL8vG4n6OfzvzRaBEj/7RI5JUAuuQXRh6Gx0WiIzQ9V1SNWXoN/lVZHvG+h0suuXUKTqNoY
3AUcOQO2vuU2WlKf7RaPxOjiDiQQI9htLdQ8BcO7REUQ+3Ph0Fuz9oGURj1vD9cY0puZ49Et0oob
KCo3xzojYErO/Kecxx0AGvWf1ZAyoYfF8NMJu85V6wLEKy74Ranzg6dgYa+FolpKdYkIeaIMoDGo
a+2bziduH9hQtEsBiWS8osgPsTabvpUdXqPsR3vh6bm5W5BOLDsaL0Z+QY4yKDTzZMnt/KJzfVQS
wLMiX9CdbxwR5jmTZXkQU5AlxPMMKRrWNI8dWrg9t1sqoDxhPUY2sBam4AUep2+luPkqJCAYC89s
StLlqWVQ5OH9C6xd4evVXPOWMf5NquuCedPNRgg0x1urc5gg/4B5TCPXdgZi7pVV1q0ZEiuh6NEz
snh8nZdU8WYdOXKoS9U7PnIXHbgYBXgQyVKx+8StTHG0yg5KB62NhPlskDo0qxJ2IBdXhdGwvL8n
cz2OCFQan2DVT3IiA+tuYjjG2Pkh5VIiuUmDrqbzn8GxaDIJ90TbCibK2kqK0qDpbaO7/sH4Njl9
83rbCVviHVnWqdqPFVSeYGmj0PhVMvr3PLNfrRYcckmUwQHjfUi0+JFoB4OrV10wl+peLyRCJuQP
mAyTdVbZwUSynP/dOZOMkFoZ1vJW4fcOiQIyEY7U62D43xCfg5RMTfvQZzIP7NZlcItexdO86p10
cEgtUTjSEBddesf/s1liQCjYnDsAq6wkf4dXkJ6qzt4elfIfhgtqArQ/2cmmEtwKv1+lEVZKwRf1
IKFYNH9BMNvZl11z6Jc1t2VubcXJ/kDrvRSdl2QbXzuvndiCzVy2g4ZBTL2qGWuQSCFMF26wkgpq
cScqeB9GYg3TSwwGANNHg5qfvtMgdToeUZIsabtq+9tsebHq1MUIOjJi3wdtgmVJKl4LwtF/9QYZ
TeccQCNKWmYHgb1yFMKS+KouWEfvMbL68vZu3r+9ic7eCpkCm52jNgu+mJkaXaKSiG3vt5qVQggn
43e5eiD3X7zZVb3C7LC5tEcBgt+13fqRdmfdRNXZFS6Xt67lGUcjb471rsGBdQYL79h0ZayWJtbg
ADLWd0bF7XOj8AK+duoLk8DyG5kzNtrqPpeXgO/1HCXWF020SNu3MEhOEvMaKPHYQep+wO18w515
A4PGkwd7iyp56qccoEb1FursFLmbztsTc2PgTCXI9SWywb7IElUTtQBPQV5pGhLlN65WzDK6Ckz0
EHFtiL2b6W/kmPiSkeCYe/TbWMLINhE0PZQXMY4jiudHPueZTcKF1twTAoJMKr9JrcB9UwHAcTuE
Gneu1XzP2fdjk1IJb1bA9uN2O+vGd5hl4GetACefs42uuKkuEIi9gzIwDE3RAlDMQWv6wa1aWGAP
II81aUeIWnVaOqeDC2IOPIRfJPOGI9WRVUVmDsndKyag4fQgGW33Rqc9Ggizgob5Scq5cYdIlThr
D02zzEkvsmbrlvZKEtBFPSxaR0lvQV9h3tILVkxyA5dGFwnMSE0goHtdmU8XkaneuNEifa9T6ICs
959eWWXlHH3BshwErt/SDxE6LVPUdWmlswBibfKyjlmEIrNjCPvZPi+LjgZxih2VzcUb6nVxw7L2
Fbsi+Iq2FZE0V9Mi6MQ+cHe4u2iW9xVlXGvPzwcQ8i48zpxiCMqc5u8mjwPa5IaE2yb/1pTqESsD
+PMFgsptxJhl0S7iavYDTRJA/I+txr33n3R7LDhKTW+gEICBG5n0f4NJ8WZt3XJxQSVt4VgMY+rJ
bKfvd0VsTSx+7zLcm0csavTU0TSp4gKVdiq2fXiwVZ2W95YQ50eBCZRdp6Th1DueavZgjlDcpFdI
VHOBUrWjH+p2Kk6dmWSvKViCWhPZya7cxZnsoMVraXElrNOmjg1pWgbCfpvdWpEMtwLJ4P4QiIAW
bsIOXfROHzPzCenz1bUWeJsgPnrBcvS0ruLQtsLXdJTh0mBG/c8KWczy259FXAJbXWtwcK/wLC3d
Cc2fMKxuzpyspC+GjhgMslOK02I7+LDr3/bs2uJVsV/2rA8dvXSw2sh9btLkxbiWH67JciofRl89
AVjO6QQw4Ks7lfAm1bd7aFqqMf/JJSKpxbrSGFuQ3MZAqLPDkYuaIzxsEQgcQCyp2majFMeiiwe9
cmJ00VDyHaLUVRiA/NmBgaMbfvuymnTvZ82oN6TzReH5qeZCuCqNsUp149zYG9nDLW2yQoghNrIz
yHtxuFs5TyVEFJPx6RmNBkxbT/XFBROjDuIr04pFFjEQXVe8PZ8kCg+tMEnSAJhTUpeJ4jlUcDDH
Oqs10bLGuy2U6g/18sDA8L0dS8FmQIPl8Wj6xsB8vjC4kM4rD+oU9bUMziBFoios8cWDfsTqJkAW
uC2EVx9kRWpfPmgT1mq8Pq9StjOcd2uKr41CyiY6J5VXYXksThByRgxQu6yN2kMz0eEab3BDiAg1
9iU3JwpSGxaN2ibrLX8DeXSOPWt3z8skzZkeLRXhN7P/J1aM2mZ8sjsPKepDJ0I+FVwN0RQ9ePCC
yOQr5sdGOzc2IpWXZCw5O9oxY4tOgjiJ/jVpAo7qcgT/ZhkuASpSzI6sq6NL+/XnBLBMqSLIXOLO
8Y3yPPevauwcUHIg5VScLQutZtL4V66V4OnXkkUZNjor1DeZuhSSmGQQqhyyUgEXOg86oH6+iez+
UZ64wpOe8p7uHd86ZA7bYDdhaurDk3Ne1ETdiIl01gEsFAnA8MazG22m/ejagNKLRE1NOXmClkUI
HzU/T3WIR3D2PFyllaAOdF7AIOqCUkVWtVpKKm6Jtw6ATXqN5Ln+xZqtf9Rl8pZbtetMmN/3uiWd
UhMkRRTlahRPbgnNsS9qflsyLNDQ6D4TeU+Dk4HWo97RGmKwjSLX1/AKmwVEE+6hFsU96/pefINh
ZmsKjyMHKCwQ5Yw4oqd7K3IEgHUdUUUKVx36IaCjoBFHhxPPB4Xsyo38hI8jGjEHW5/AfWnYN+zR
Cuw73B4f9cf7Yc2/B9EhdhZo75nbYvkdSkIHdpNUarWx/Z8ELfqNuM2+/+4hUkChYURoIxpcIfYh
kQLAz4CnMtnSLBsXvElL5iZTCDnDv7RFgQNAT8kYxeni+pgdlO/2d8sO7sCWLTzDqYD3KyvbeNM3
EyRp4qxHert9QdI3JL5MAsZ3GNVbB1aJtStmk/VmpJsZU2/wC6xVwuKNU4npgF/nf6uWRhPXhaHs
ekSICJHg5qo6oJNWRSdbHZtUSje1gLjg+jnriXaXOq3LO66oVfgzIUQCvm+wB1caSk4wDzq6OM9e
KnYEzzmnudzyZeGLGSWm1DExRA4AfHqXfRcWZFLmC9o77QP4Z1I1P0SahTCsrmNN3eqIKxcr0beg
5Mcax7VcIWWCJwTFrK7miyLdaiEez707b6VsrySanaoq4CW7UUNVdmbLYoKZv2a2+iGRL1GgTaFz
QXDHYKhmllGPsGXOVqfjvjkR2tyq+vchG+bgE6QiBoY+xwNlrMUE4TWaVQpoCK+aYIn1nLMKMg/8
6M5NkStdiENLM3ftayo17w3Lf06fzuU6d8niO9EYvk4yM4FKutiaqWW4J9i6JzghdXlHg9uh9Lm9
DFRAQWviaqW0hOtGW29psuXTrI3rIDVejWna+lOzM3iKb+JJukVSiM1Ojv1YJJZu50bsQ9rli9gw
dscyWTbb5KkcKzZ47sUR6S6CRh1bXV6NDDB9mZ1dziONBDmbrzFRfHnrDb7C/bB0cjYIPUjkWUQf
L488uMpj0Av5OY+JIcM0KFHPuiMSLOmqiSHIZuCTUVnL9a1I45y6LChygYFi1rSJZRmsrYyYehLW
iGnK6J7JRyUfrXL0JJbYv19ygju/1kClyfyyyAJFDhQcxjEuHutZ1xCdAnJP9U3VX905dqwPy7+F
2Y/TVZa6WtkF71vuDYa5/V70HVOJkT9esjfKQiYlVS6A8/XqzuCtGXhhG5D8Uzajb54LEWK6BL9+
NBiyFSSdAUSj9jVYdR70TM38Hv23eunnVonCMltAdgBJ95DdDSibowcyWrOabpiBV0Yf59rzibaz
EwD/UD3RSLmrbLXWLog6KUyjOGvTnHwilFcsssh+19++BosF2J77DtJ6iqh3pPzFZIVPCIHp+kue
eIdrBl5mbiKAHzgZYRlhwtb+6+yKDFrNqQzVgmZ1lrN3gG4Ej+SxXxe3U2iZIINlYjMfrZyy0aJf
17XZ4zYYmLF1Svj4kyW5SOPLuB+M6ESmLDkaOFHWH0QSNrWQ+5JFrSlJARSxjW1AdwqHBO2Q1zK5
sKT/n5hsUfN7hFhlbGYztb8wCbYOAy2tO5/+HOSBX+f0I1ckG4xgFMY9eCamP4RviV/E3xOR3+s6
pXOa4Dbc/8CY0/MpwMbeC06Mb3NsMxpSDJi6L269QVXBL+t60NX+0OpdhyW1jlkLZSjxBtWKUlIM
mFVisctL0z/3kWbpXfNdySbr+F0XqOrosRS+LV8X/Cz1upB2AFya2lMkVhiS6teMYOHpoIa7eZ5d
N7FR9llneMql4gRWf4jrfEcnqps+QwiYUACVJ6Cg6D9XLlgqpNDgtLL2J7Divs1yAErwc2rMgnZm
ZHZhPO7QRiGpHB9hK4rrlR7RLlAFKL41SZRZVri2iV4lA5yrU7bDV18M0chu8tD3IxO2/UAHUrJ+
8ZVS1gpMAPB6MeOcAHgr0+PeebEWo7RU0VASnjJ+pzIluEZ6BxiH+SuXrEJeKCZE9woNlGkKXN8U
drhYsqwAI+MtXuBk6toh/fdGjN32HF4zMHRNZzWBs6ntrU7kpmLdp/qwa7iOQGMLcbQTmXQ/Ig4R
d2PBA3kinqYF+fqd/ZktFavdzAoJ6YY6MygxpJbH8U4mXLE/oLV4wG35t5FlNn8ag2M5ulDKGVye
VWeoXS/4wj+WILNRApH15FqyqRTm2u3GQyfZVSnUWPeOI0ZRul6uU++FbYUJbvsNyAPNeLH9b9xd
4qEIEPhqRi2DmC7n29sPVxD9dkTp2d0ohl3kBpB13ln1v/dnw26y6JZqFdc/i409dVNpxlz96AFs
GndnL2fIZ2GIZFsYg4WtXsiz7gPrxd+gwlinwQv0abepZKYXKY7YCAELRv9OgyUBQwKFaNi8P/KB
kVNFQU7CD7a9WAW9Y+0DoJOGrOUaltzEfDR155qgSIow4ybgyDkTlw5RQmjseQek0H9ueopwhrFt
F1BctIxU1giFr/z0Z2L6++DCT+o+RU4ls4rh2jBFiumCEBvRrSj9cK/0ERrVOeDgJ1BfqTw7woKe
yzuSqbhpAhJxtOosuDQSfxMq5/MnhmdmgZtti6TZfYpy/PkOP26FFqrjT/OkDjolR9SMHfyZ2+Qa
wQMMSOvqdKmT03/JM4/dyPR9YazLjf/zs+Zhmexy9fHiAco4GmSx0oCXJE+9esGcChYR44aGuWP0
Fl5i6JzcPHwsTwfMvZSOIFRxwZn9iVBsIW/jSGeZ9WTeoLl/Z0JF2SrGem/jqgmDzam6VINdp7yN
TmLdBNGk2at/gafCw9FQTkmT7nB7bbMUVvTCp/LrUIREPpnWzqWc7KCRaocVF+JY8NKE743pY5dc
LFz1D+EgffmpU6neWgs/q2Up5MO9hoacjOz1knn1Tj5dpijqTjDldQE5Z5MS9yDpQ/SPjOqd6QcO
ojrgKC6V/v5sWUi2IFCX8IvjYSEn2uTprU0ySuUUVDvxkqKAXZKuUdN/1pjNuN03vJ03oGS1nsSi
8W/qxx2+tOMiRCJfta34N0gY1eDSmLXVWDhnlONQAWbjyfMnIz0pBulBll+D9k4gryzI2ZHnyGBZ
nz/YVkv+yTbnfoZSGEy9r4Zo02TIfMlqX+0inur8KiVoW1VOUh4TyHFvFvzZbyxXvIX5SpN+J8Pe
gC+4jAe04oozxr2ExCo3Igwh3DfA7ZxS9opAM/4382lXHH+ri/IV7oj14V3sQsGxizhCkGgW10iB
pWzTsiYFQJuBLzBAqqE+IPYfVYERd8Qu/4yPtEf/f4VinQZ6bQ/Vst8E4GeeYekYh+GeBQZqcC0R
Y15wnNlGDcL2E4IzkejeGI+dYRXGU2sfxKrPrrVHJeIlfiGvRF1/C6W8mu0lqA9vxRE/2uQqIJoq
pBCEQRNutMSxAO/FSRR05IHf+oUQWyhsbsc5dvnJilrF/IVwoVD4hXWQSwxdfbfHn3yxBiOIOIgy
6vfotOPnUuw6kiPHh3ZgTDugOP7dO3xLkdPaVGYFDYjP97+wTfjV4KkH3GLXYyXuXoT2XmpLNVNi
ymY7/KXkSw0BB5HXoZb08A57vlXgvGWToHPxz03LLJZFlu/LSvAJM5DQiFGrS0UgHlXwKBvMsFMr
BtI1q8qAbKXJNG/n/5HBABCA5M/LVQEEuyWPGeGGdxaauW6XYj8iLlvb0Qqm+8r8pPuHVs970NHF
7SeZJOzZHkvH6ImTYkvZad19QXN71EKX+lXEeykt2Jz4Ina8YnHxV1o33cYB50lLYPTElwpwHPUg
liFe3scocOyWL6FwZZKaPvOadenrmGMpa+DLpPvVbnCA9xagbOpUvRv5+peIYivyPyHFclB9SrS3
/UyVVF4LmsjWLuqKB6F45G2lU2UcV7brxnmnB2Xd/i1xUK0GQT4IX419W+rvYYPsSAt42DPg+C2b
FjC7ehF2SRp686Kkq9PvRaXFgqM2QUQ2ssU15mYIuWUt2VEzY898Qw5ochpHYcuhnLjwWrZhGug9
oyriPLeWd2wzbc60ZcksrIugI65TUGM6JBGYS858TkpW4tnk4YEz8Pmw0Zvlv2OguYwB4fANisWt
AnLQFXszNQqH7Sl1Y7uZ/XcdHOvl0hDY8xl6uoA00U8IDTHB+jEqt2l25VCYVrN8qFCF1sWITvgN
s4cGuzA6Kd6HzVKVKqCOrdntxHGhmVm5pObzDgusOYN/R6oEsUkomU+N2+mOSiWoBI398f9lOWcj
I6QQxuqNigcv5x9gECVhvr93woV4QM1KnGyR9wi55VLMddWm0OtMcN9YGJYcfK1+7L4PTgXWpE7a
qIjT1+7zt+lLoX6vvwiEIsp0+HCFGDiyG4z4Vy95xXVdyI97N7aF04pNGcfmijejz3eli11UhDaf
VViI/fW4Cal6Nz5IilXiizsl+XYxdD69xT30qufQQnVHv0UoSMy0OjC2923Ytofb4GjckGT/TFhG
XzZcZ6k+fThvMKe+od/7A6oe2zsjX3wRZ7YnMjY5T5l7Lu+eJiCqjBl6YDKVVFFwL8qsLRNcJF6X
cgleTSzxeGCTpzRH/Bho6Rqm90qhN5vVWPSFzmVBMq6yYLxthbka+DXBuMhfunp0ow4bTU9f++Ov
78uJdzWJ22U8OKxd7B0JQwbCU8xBncBQgbI4mVmY7VHyGy7PucwcJMdln7RNxddFUtCWzY5XPmXw
LRGS3LyKBXXO3ivA6uCE+Cz8LwL2/9DvV/GBUfsaZPwGWzZ+JRWzwum9vcRtWTjHQrJOILuqVpyb
0lWJYsM41MU+wjU3SNu7oXN5BNaB7tseunarE6jbK9dsi+aecVmnLsMaDxcPuHE4cbxgHGRIK6EA
SGKz7swSmX+f7/VQzloRxEL6OB0LflhvUxRf5nB5KYr7MF3y2sCZAAFZ5ySW43GyQz0/FVL8Ogc2
+GozKwLo+haKrm7Ea1fFoTssIwDpGaodolU5z+F9rXPZVDMvLYNnMWxqIejtqXdfKe4V+Zf7mTOn
iEbQC/d9HAV89/xDlQFEDoTFEROWBCxCGkqcy/ChJoiDH4kcPe3syq305HVcsGt4qevcv6dp+9pG
wwgya+yznfWTR4sZRQpl1lXD6MoT/h1NRRnTGgMv39NOMBGINlV8WxitiG2RTJZj7DmYqNQXLIue
Oy8r+TF1LqCcxuuB9C0kSYIg9qDdDJdfWwMzD2Pg1tcedTTtWvFwUwMrhnWt2LHmuM+PJCrodrpR
E+pvsgYZ+7Lb0OpvEWkffZM1yZ0W7ogjrEws6fNZwIsO6M0LtcLmwuBck+4QktUuRStm+fGVzs5E
AfUZGXlplvtIfsTzS5XVdYdej1YhYZq7nDCGVYUkfScH4MGEXrBSLz3cAyBQwpn4Kr7DffvRvvDf
ErfyLPLD5AIWwD/1RZA4qB6p78mQFH05X3+LFEeRt5txatzXaynvSaeqEhU2QvY+9yDrYmmlBzgL
KGcNCzn6NGpI2MrycY3+C+IF6YRqCuBg1qaokKgg/O3RmMDliDo9nqL0Tjjo5NWSq8ywxEf8aC70
rw+V4Yi3uL6/M+eHMxLZBYS0Bl5cDvMkOZYw31LLc8zur2kBGeb7etF301K0v9jps9r0uNTa+MR6
cbgEvf6c+imlH1Hixztg7OFTYAUtYOLtMcAEDxtzpa4mK8+AF7fv2L0hvCk6II0LQD46yR2CI5ji
n4MdiqUZMlHqWX0JAgPgKQGrZUR/J99p729DSUj97rbpSHaPmvCDVjmD6sKCIleaQbadGVQyhx2M
kv8pmGd6qNKmIpPUu7OC8OVgUMrCov1oJe5ky7AC1PTAVnF3DmfWxp0C6pnJYcr1iCdC8B3sCqUk
LuGR1N2hFGEbcBJvi6b+D9L3qLNpmlxyIceZDNNV2u9mNFGMKodtG4Scaug7SVNIKqUqg0wQfPqR
YJp2RF29I3XpjXvLy2G5pieUtaSuCXXIut1UYteYeO1Vu6U8xLOGLVBAzcSW4r+ysqvi4A84xeBw
ToB8mXs1/0uMDLxUtpY8jcaIoaLR07YYS7Xjk2wlpjcJZigqQX6VXUwWp/92KznfgHjNaTbXmeOg
d0UUaSEmmAA56Tbp137dkWWcTz9svIpa+qGGvsE4BzjGnfF3jYaR9O4uBdzvXTlespGINt/vYpmF
pZsMf204tKing6D10u9Kn6HnKo+SsaavsQ2rGZ1zGd6tgf58bGsQakHrmeQ7ZZTfXhNeeM69tjev
FI+aMrSmkhc5kwI5CM9EaBuUQ6pX1dLwqes7MHWqotL/DAgTtbmuNjpqfhqsnYzWbDwXPei0tTOI
nAkrtu7ErClt+ojx1q+09AHKyJ6qRMAHXcnD/z9v5Iv7ixwe1+PqKadiCPooRl66XMTjA5ENuNkl
AaRvua/ayNnpv5je0UunpvJGKgJLd7Z+FGv8DDXqvlilFms0o+Y1+9AHeVXaeJx2jvl1h5Mo/HeG
vNEMAKPaJ0wZtQe4wJqLnnfnyR7evZoIX1vfDX+tOR4BTvv4I0vcNmntFUgfw0WUgUm6kIDVt8hv
z5lB8hyO432bNvy/zuoG1U1l3t8WhRQ/YlmDbC68Q9ygWHOfENHmG45ERMV71Un/qcw3bCNXoUOc
k9vdNnJ7I7qwZWDCRkchUGFgwsSfGn7JA3Dr40arW8C8uhy52avvWgGT64sP8bE3o7ZqJZTXaTUU
YfxU9sVhRtBfUlbHd9DRpXGkFwfbH0htXSrkxmVMCrvV1m8ZO/emo2JwxIL2fFgEAMY1F75hYQ4I
vrrUIIDaH6p/Kop6UZCvL0o+NHxjE6Fd5VtgwDiGfI8J2p/cBUX+BaQHOYUyFwFO6LawA6sujQpz
QD+l2NW2ghAf9g3qlJA72kRnn+mYk+IzB9w/5yWIv8+CDgZMRqTGyg0HMq0Y1OID4g2pop48RMjA
OjOmNYRUB7wdequam4jkTr6/mJCjzZ/P90ZaYwaCGLNKsKs7x9QK54M3M7TRq66OI8Wa+DdZJIe5
zAK/xgaTt6dYFXryUD/lE1h6r461s8OCiEQj+IyG1pLX+ng/zBLMlZlSp4P+0uBMkxGv2/iITh0H
pNiYU2wk/NMzMhAu+nSJ+3reIz3NZduDdCXmSJ1hup+JRRG3qQAo8vOyjxaUvt5PNNiPWYSKKR3T
/sS+VlnRDkMQ2k6GyTRUVhzvP6Bl6fiOlZS+zYwLTTc4A40YPpvReb54E1G2u6KxvSSw4fNJyrEe
+XBZPK93cA9IIjQrRssxXG2PDZ1hxv+d2UQAn1o2uEvDRzL+ujbw2E1nx9GVubXt/1M7UpiphPWz
F6o1SqtdewKbZVvKAXWDXG3ONlcouhURtdyqjZAQOQFAJDJVoJwZRdneS7BOIlnj0VgdWg8NaaWj
oQMP7g/fexxLjhJXA1i5SyIdAxbvgCJhbFbqezRLmFbnCZKnOLZiIGNpNfMReTCjTsSzG/DZIK5v
re+UeTDg6Eg0ihgxzWOnYq3upVbzUP0u+E8Ha8iIS+he75VkDM+X+Ir5TTnaZ4v7m9j+vObDUvsD
+pD5YlwIsAk25uBqJMzOgyeHOVmk5yE1LY4nLs5T2nfQFTCz0aYNTHw5VlWsyBwHSQLzDOUangsp
0FqUJ4W3YGRJ25a7XhIVrkNbBouUzZKFMuW2xl+Yg7xK3H5sohqJXSdcCYZKUpA0WoXe3X6MnJwz
jem6BpwxUJg8M9vYTjyfeINBjyOl1Mu5FISHWcAr8DyAibET5C1ZuekWKygUzkUiwSGkwfksNK9I
Yw+dCZMI+OcTbR31OAKjYLXU9phNJU6/SGtjHfjbKWxAcAnxt8aRJIu9pVBgSvAQ/L3gzKUgoiQa
e4Qwo4K0zJgxk+9PKqvWTYAupMfo0HoLagC3chzjVV5T2HExrZVUSlHrq76Hxy0eExHKQv59XQqF
ZkzSwheCFEMjS8NNbh7u7NOBFypZo4pIKmBmMnP9how2fctOSA6aiihdmB0nj6QkpKYRuOcWISga
sF/Zk/IgTauaXODwNNMwzwwExen12TSJlR1YQk4cCzzZdU1Rpg7b1G4b88mxC9AHOWJvosuvSgr7
zaFR40lEz3ULJZxXJSmKQqy0Z4lRpCgCA2+8X6otDS6Bcg9JsEi9/4j7Ebzu4PVVGCad96kFWAPi
M5+VViuOjB5Su8P4EjlNRoAGi+jQuTdy63NryFb/HqHuTRXz4j1c6D3tv6Oeg/G+OThMeqTdEzId
ZiykUswPRfv3Va6WeOKsUoJg5z6PBtnRvR7C6bquzGPoeLSKAoVgEpvLUCyoNr61OYy4TusoY5f/
N3ZlV7BZf2BXgnxnYnVXaVWhuNRS40bTtoWDlTlA2JVVpAFbueYC7Zm3YZfT0cr/DVIv6rAe07NI
A9Jfm8u3Qezye0SaBSHGuW+BoRzLQK7X5WMU+p2hWyxAjGsU66ox0PpE6WKtGS1nVYJqMZSpdUmx
JApG0AM9ksaZORDs1QG9yBc0vMeo28fL1n5ZR7gEDICuZrMl78tgnQ5rpPPiB9AEkGVwOyIhUbEd
SkY3UEuEDaRvfFDC3CCK3d6GGgW5NRRN18j2DtdS0pizCn8Bg2jhUY6dSL0W7kGlSQ6biqK57LNc
fzNUv406Q9/laqm1YZMWv3zXkIpOx6zxQcjakZUpo3Y4jrx5ua9I6qJnTrwj5yuHBraY6zVRocW8
IbXHqwk2N7YuSNlTUl1cH+M0AZGMU4w3RQXm0ATNhhNsgATddJj72EcuDZ5oyN7Miy7MCwUtHUPU
vG7Iz02fLL/CFMjGV2nV0YQ5DlH0xNuZ/rrFUCtKt/A6MSdGbcR/lLjgxNoQDnfJH7Klb3+yhGxc
Nt8u4TqADMNUd+VIXIAs8vMdmoqnePl65SvXQ5z9OgX3bYAwirZyNBPqVFSZczMcHZLcZlyacL4l
aKAT9Ei3hHqoq8mCxfxh6Ux8iWWB3nPae+sz2x4C9XnQNa2CSC8+gPN9G+i8A97dUyL7P2as1ZBt
QsBJfPT1F9vUCGWNj8Pc2SWk8qAuA9tgn8nnIvqkPRlvlOuKh2RsBdrYZUzgAPgcaQM0QqN0Rogg
7tylixJr87joagr8D0duflyDhVVl+6H4l0zfmVgOMfBRd/RRMyDPWfxiy2k3ra6y/0R215kjmKDj
esMMCsydKbsmBtLYO71RYPiGlfv7kCihilhDmL5QEPzqRIVncc/WxuSUJSggPrdzvr2K+tN8KGVP
4jvZvvMTCdydsaxbaIxmoDvLNO2YivKbtCoS8sRJOIztVdVd8ccZ6JQhjlV7xM1kFU44M5kqgXRw
lMWbEosXs/+SetFoC19Nm9jjI0dKA3HDRpIL54q7yM7CJkqyd/sARnfY/z3heYDOrrpX9gFdgVQk
jibip90FxfKIz2QTxaq9myjo4t5Yvmv4afZud/s3dm/l21fNosGxMvfAYpC9EA7Z2btwf9dExuR5
tWGjooqubiI9LLkDzgi1bN0uCbvOV5LX2hIqvppCEG8hJai7i+Wp7PVwCy3AV+rImAFlNrX/Dgf/
LHEaZurw0PYQ+cqMy5aPR70Is1Nv/nNU67Yd+vac3aVHmKqXvggmlQtWJChid5fHhcrj31P9W07k
jWDLE+RBop3Q/mlPGcKZtlMjfO6xSckWsNw/9z+BP7OYHjgf8vicNTuGIHnXfoFDQ2sbIHsJJgBU
3yqVc1ayANQRFYrw3T+Cn3vemIS0kSmbO30rpAMzcCxBFqNvXdLTn3nnLNnWDHwg41EbWLu4jHKY
f722ZoElYbgVct53RTyZEvYdYJnxYNyMic8UYDfWrtXKSrCWL6kh59YnGJDKF3LhLB2w6/90G8aQ
LnRCU5I/GTkuqZ/fPaODwcWrr9bvgEK5+7LY75FSkn24+M88VG/McyDnosqKYAGkMwc8o6IN+zxE
tVrtKaLvysyFlKrD4ayweUv0zoxHepGCZG3r5eFEyqTB0UyuhNSJ1VfZLkOhQwLWYs3105CGJnlF
TwfaoK1CmqyQGiU8Fj4MOUbY4ZLTmN+UwHwxhZc31svoI/XEN/xNoqqsCUyPAICyzllkIH3aXEQj
HBlto40W7RJ7dzIeVNVXAu/m0en8Fps85AgRKm4syNpHLTSwxT8uvubBWZ5GvQXrqOngaLocEu3n
iNjO1mT6zfXspdqCFMki1gw2hIAFFLi2gs2YWPxsf1x3o1af8crYg/jfkDky6tyvbXZeWWL5xpwI
85vtg/DXc+/PJHVBaNjXtn+FjBPL0CIi4jsHQsFeAmSEfy5gqSAHqqjNcw2X4/nuqBYRfrvrff+b
oWS+6fabZIkDYcmaqycRpNLfMS1L88CSY3bEu2FZIfQlqfRWKtzF+J610hGZGff/nr0u8bKRXsGA
bd5no8Ds2HEjL4Ksk6ZO2i/OjkVyI8wjJypmR3QxeMGwJFC4MQNvvFtiJUKsadlSmmdaCK01Rj6O
YVIENLNN2m466XAfT9dWtz9nsOMz/E4jQzKnN2tNEJY/nQoazxcL9KFp/7pzelQzTZN2aRaJg+xd
qrzOtS/0FtA5hheQYCm4p71rnD9bD6bmbbl6hKKeV1ZJrKp+z5FlIP1p8y3dN8gejYh250+zPIJe
9c5vs/JNkxIJcHBW4z4wpzequhjXAqZJf0BkjIckDl4bcK+XI7hMoMRoTswVLhkzMagc7HmtNgmL
ygWJJjXfmoTPYPf8teqNdibefkaMIzw/4nvOTSprgzKxbsSYP6T8yUe93FAAvIiR0C0/h/K4U/B3
pvJOyho0PM3otFZqG3PpqGIXIiIRhJB8oJGTpYpCX1EewTwgTJsOOC9slwXttegyLvAJiLQUXPTp
NFAiKLB/6s5nntal8MuP8G6NKIrk3/8zou1jbx4oJebClcUS7kw8OkqChNssP/AMa4RxDCyXt71y
YVeow4CkiIh4P7BHxzLG9PeN9g2ANIoaoWv1e8ziEpu6gR1TazXrqO9vTefOpv3C3B/kiB18uzFf
I45hHDmTv6ZNOVDGIDTSXsSu+W8p7im7KaShuyy212nQoUmUXZfXgunPWMzPXL2g+bamZmjdmtpl
rI9M1SQyCpda+uhWDtD6NPbNTjTZsMRwxih3DLyuf+aRw1u0pw+fDNiF0Ipog7QVrDM1i5w6soVS
mt58u/WLf3tNesBtC1lP4/WXXiyVVp+jJ868dcPM77B5VOkhBhgNn1Bi9cvY+3b38lqpfcj/B+//
VFDPupmQjvb+FPzDv6b4Lpsj6OrBN3tWFxAepvWHx4Nx9aIqDxnIl7KSTeTPLDXZdJepD7+tieF0
MFHMPu5pI6P/mj1aE6TVKsBRCH30OvwIrWqFvM5cnoXTcRzzQjjM4Z+Q4Eowzl5DddnnUlqRTvO+
9nh4AIxGuJs1xOYnrZLIUHvZpTdWVVt4Chs/ZUc8WS03B4UZW9ZAd3EEmRwNoJ9MaW4oabyq/PIX
03F16Cil05PjYsYF5ECQMfqR0jpdPmeUsjLHZu7ndmwCfv2m6sIwI6dLHFpKE02sTDWl3IRGD5Ug
FFNivBcMAzk4OsrGToD1A1gYIfToJcxL/VYXRKR0pbWZqj59AOuzWa0zKddPnbHYV4p3St1pjxyl
7By8N1+p4ttSM9cHyqIG80ifRSOzqRao6qrB+p2FvHTufJaQ/3iPCYCNEPXOkRNpEXT/XKZ+JHwe
2fEbXHXGl7K7wDulw25NaKkXP/fLj8603IXnTQYfEeQnrhg/+ijM9Jq5XxR6WqX0ocUXVgUH1+DJ
nkEuN7xSLB6NuVwrh7bIKBpvcfcMIVEV/N4Y4Bsynt2T30q18HBfJGeynCijzHmSh/oFmSuF5QJp
3PxRs53BMAk2jKkhOmah916ddjqfa+DVntFoBtHEQL83Qaegom2uiLHln5ixU90ywQEgGG8+UtoH
Z/CW549OFcnlDscKi8fWev0Fg2bkf8TxvDRp/co9ysACouNu+JYlh2VktkCKLtakNRsLBsgJ1K5Z
0Tq2bEJKvIl8oOMpHqEKQgn82s5W+uR9gr7f/NxuxiSMRA9nO26RUiJk9Db46aW75oT2gzA8e2xG
XfORuNH3krr2vaVEwzRj+3Fd5d5eTUWRQrlwxVmBdYU6rV9mhwOkr/OG9KR7BIIINtb2fN1TAynT
ciFsK+VPy7BL7yt4z1xMqv3AhH65+dC30Xh//eaw1sPepvWFHdiMV8dGVo63xMSQW/nswY9oENqT
DvipflRbCUk/mL28lR2JMhfSoAZsWSjauEgX43hBO72vWMAKPjist0IzkfKIP1Df8lG28putBSHs
GnVqZIBspJQe1045wz4If5zumZFKvQxiVD9R2a+iPZkEdvDYxtfps2ryMwsWSnGZtmATae3LteFP
o3aUmPS8PyrqMJqV1MQwIA1wwC94yIISP7Giu6a3KpIw4hc3XYaqqyEg3KIFCPU0w06Clh/oZUtB
X7jnBprMsawWQd9+o1VWkBNKd3XaXUxgqmSzbXYFS5OPrLlcWLSH8+X5maWt6yiwqEQPdajaF1T2
XUS+mX/SFeDf9yE6+UBw7UX1bPa3X4OgQhiZh+ZV3yLDXJQzDeuX8nxdqRcZ+8naz5SGJE7Cmsef
FVHl5FLhjmNNyTEmsaLmTp175ryaW7FFEDJsdgxe3IfgvflUjka+hkuPFVW+hNY3kFQ3Oq0gNv2i
Y0wgDhUpeJKsk36/muFJ+7BLgX4CnLSa1+awUJ/JXXN6tTLY18dCaTxuIp2ZUyAQN+C7fOmv2iCA
ike+x9G3I9ju1xScWktb7vGsGw+G+XbY99PJPz0fnb+Ws6wD1csDvANse3cDSNkHCY9n3tt2JMwJ
+16/znQbNNhR0RRtFybPWI125j2We/1IT9CrQY5XApnDt9YBdgUxq8mhwgtdSoO8OOPOpTCXEWCr
1Ot6/nPssYbRJN/LvSWb/qutfiddU1YhD3bqOSVBc1kbyJq6bKOVPzrRoOamz0bWZpE4G/Pm5Fkn
17vgiStxmSXzwAt96ngL386SR6Isw/dr9U6nf0T8Kc8bSEkzuyfgVDmqgT7ZkBPLUpPi9x4tXjWa
sgAOkIPFGA/A/49BCgYPzaSwVqbCpaESsCml0a6Cw3bBwYuXDhpwegcIm61mV0CUddjdD5Bpclwu
AjuT4W503qMJ5fL/mVAjnYGkicVuI70ZqMBwQSWlr4KKB+5NurIAJnH64nIZXu1ROlWqNQABRjh0
Qgwoki6V7gHpSrxr85AjyiHrevLPCW+IMmoeiTAEhlliYDBdzcmWNXdiy4ljXaKVbLewh6eaRSMl
1DatrmBJmVCSlYUPsYmdy/Vdy01oz9dPmJ+XCRvjD/ENSinF2NZh3lMGf/46Lf89/M0opZ5o8VGs
lZDIPfwb7e/QvVu+I5InY9IVNJBb8p/bplVAIK3kdhRZcuWCTlHl2tEATxxHKXWn8UDTAv9k/tWk
CtWFa076y5FUCjbQLs+FT/RZnVrZEFGMTXZavdEjap2nP/BEn6Q3nenB37Ho3WsYU2ZtlQhj7DU7
QbZ9RJG30oI0cEviIyhFhqUlHcVUd0ELIG2Xu/SZoZbiGojR8y3SINC4AbIU/whyy4jeYlkB9WR2
yo/ZiXEvnF3h2fQsZZ807rjIjJwxDKEST/LKJ6nDF1cv8kOhdN/k/IyPXwUhAqFiEEDZOx9vMTF1
7TgFs07NEJpEc8VkOAVLeFH+F/7s0ZtC4NVyXY6PiXwh4SVEhfByORm3yK07X+vZUasRB14xZO1U
jWr5J2j8YDLRpKrBjSDlDDbuM+tUjgiOatjKYud6GVstgeGi08Iaf8b/FLEBfX9/G6j8Pz6tHtrT
PrLjc3d/HZ4COI6feGQD51pNRw4dX8lNlJ0ONHJgFkz8/3kUOWlC+oGw5G06Uy1uHqSXhKScF3Xx
C4xt4zQ/i4P635b4AZtKm7EaPciDRYKBC2/dBKna27ZNhu90uuGMgn/cSyGIJFTZLt8C0lRRNG4t
Ciql/mhs2UWhboz49GqpV6zWo8R0iYsAZRMqUusVevkylutjPV+CMMHyNsEwrHgmzb3nqq54Ep4A
283mIqAx/g6ViZU6UYXkUd/BVIbRwi3IWc2Wdqy+uu/F6HBReTymYVH0JpD0w+awVzgdorhz90gE
hXALoaZqu12CFvcht2xL69GcgVlYIeSau7X3mkmR5az0tHjwT8dRUyxnhvS6Xqjm7Hzge+ACca3o
C6728cborVtOB96omMq3NbjGfGmODwlwvSSTJf+2LjNZeoZDvx9eBhNg/kKnsr6nlLBOb5nY3tOK
4rDFB2pXa5Ox/CcrCbtb0RUKQwHuCmojEuwL5X8hh/01hx/hMgfuzrMQEtCx96Br36VbWOVPn2U0
SMUAqFtGoN1mm5tBp2yp38/zbq7kMEB2KOgGCN+7ull7rbLe57JkAwb0+R3U8GotRCZDeTrWacGZ
METm1lHQVAXywAAIskm9lUGbmZR5U3/XkkVAAsPyZIWFszQ4nPuRXVxOfA/wnZwXhdkjHcZTxSyr
OD92w9bh9fJDUfDR6K2wkmbJtjINSfyehnPog2alB3rFTyVxPliMbmIxKcqo7YxRssO9i4juaZbk
9HvKdA95X8IR/7lP9C09mGpyYi/ffv3c/lrq8vFUG8DgoFlMABUO7/0O8ggQjlcva33mkCStjxg9
E+Z65WVRCDflyKyn7jBYJY5LU6FuQ64kPgnxzMEEGizObelmmT16omho6dA6AoSkquDlHrDWRn1D
c5ChLvR3EhrsB09gsKiG5RxWoTbbFTwVI6NcIlQfa9FVeH1Ne9O01OAsJ1/fc0ItX0VyuQXnSSmh
rhQCKGdF8z/ZMN/SNfRtoN208Hwj3KZbOU8RHoBOA4QjNajNhm1l3UdNyVvtxdz58edWEcnhGa0s
xTfT2+XocEV2LgG9VuzriKQBS0cwO8YzJ8Nm1yXzIMOsISq5uJ5sK/W8PtHlJGb+zarl0rnQU9d0
dMbRs4W4uNi6QyIpKrX0XMRdor2gvYh1CBTOfMndKxyo0Lvltgf32mBYcxbd61V3xorWDe2hwCKS
hkMPrWO3tp34pGtf5rkh79Q6XtZ0EYO/54KaWOqNnezwEjzIfpameJVXKi8rdiRaFO03PwD31fHf
2uz0vRN1Zj8E1Xq6dJDJKyWiZ/qj75cWhwBTjLh4YQ7xRHpsY+XOS6MusgPCHAD2goRpHLdE21e4
4KbMlrIdOJL/pamthb5gYwA1FV+qOsh23v5ctLf4xeGyMXdhqMNtL4B05O0W1zUO8cZ84V0lYJVd
V0ujk1Iv1swL/96N5tcXTz28ax54pv8qfkVFWINFcDbXzziohm/kawbhct8wq+lxVrUYFWBPxdlC
Cez+nZ02KNu4oiyPPg9hpaBc0n1pTYMitQcLTpnoRZplLxxcz8YrIO0t9v2SiOzVD8pAiDArl3mY
/RzbPQout3mm6YGnUph6GlJqfIlNZOa8E7qtnsAG+etOMdwdj9i1AfKsZsQUArXaxTw3ab6NAdFV
RMarulUgdo0SZjra8XXAvzkb6PURDw3jv2/BziV1wgvb8Kus9b5ulCOoHvKj39xA5S9CXwRNoqK/
IJz8Wjj/XHgvnCfBFRQ1TaHrTrbJzVIZgSZ0TSijW/SELLDphiX+mgwwLTATeEvGRQZsup/ZgHOd
0Ia0sS09lseNf6s+phiJIhi2KmkmJG9e8HLhIQhRB773Oe/fe0Jl84nHuzk/EHZSLN6/Lyr7AWTt
Fp2fiY/A7Nha0vi6b0qairoqQgYYWxpUJBM0cGhIsolGZ3ZtaWg2ApiIMDlr5WHI0x/SL8FH0i7A
19io8UVqeUw0e6UOJ6FBy6LouPmJ1vk2+5qLqp6MJGe7xnbJEKbX7J4ZSlu0NTnFMtWYYLV6banO
rp4pDIsTjI23LE+n9kBrQW6Op6Kul3gWKiMaJOBT8Pf1A7+VLKy/ZHGjhEsaXm354Hssk6wCw/YH
gPOs8En6eae1I6vaCQAdoHyiPb9ux0/j6vytT4wQcm4SOKPYUokjTKIlHMPc4xcL9ZNBp87y6HY7
3PbLpq5ez+8jB3EEPTQvyIm2zIBCnWYm8VqsuuLhWS8UGLwg04UrI99CPtayly/V5JfsRtXOBd0Q
gbRC7qPIojLv29h6xVKYmbJVbSeME8a/BcX/fEizvmJaQw2naWDsJJBDuB6osL7X5Qs5Ulle/1kv
wqPw3ZJY+EvQNt5kwKXBks4ssEHUFbzRvicRxNpy/ok8wfg7nkfo1ziDbvQ+gvqQsGhuq5sMWzQp
SBD9YNvufGVFj4Gr+32aFMVp3F6O3dRf1nrQzMbzNFEPVn3h4U/K3yrOzSWOnsDCYoPcGVWN5rIx
nIZuudEPNmtCM3LMmbQmlbH7aPBuJ0ZCgybsUe77Yzb6uFJBl68w+ET6D2koWOgDCK+lt7S5xIbo
oCQcm97pfo0nVgA+5yM19PUCErOXlad/+ISZeln6T9P/fon6BN1QhGTHR6kRBi2kzUBJiunqBifT
QSCQ/xgpneOQtvtLe53EzZJXcKPr1VOl4+OV4xzhqHtRfIRQ3TxfWNZ4CjhPWNUrh6PIBiOiQBrO
//fA0Ed3F3og5jIsRNDw80i4v7wVVjmitMZDuhhHcfceKz0xTS5kYE/YI6IOK3eT3D6j6vaqcNuT
grS8fBEYkmtKpiIoGFjfSnMqA0KxRqzjkac7PL6ybZyhVQ9GDeUnL5BfQ6157RpuLKYwvwJVNBX0
p94JG2E1ipvuVAu0YCoy8GF1/OGeEVTyR9KwL3qyYGQ4sQoWklayUb2h8s0Age/kbrMPJJ32I7ig
kOYlzzwRi9uzRQE7S+L+HrRW9h/P2+duatlAxrGub1hFwm5qKpyyYSHr5ClmrNaxVswFXPaifL4f
KnfxCvNlgzV5L43Bo593RWmnZ6ZEyJQh7scHalzFvxagFDTJI7rIXngXwU6qqZP+qLZGKFndF3v4
jYIkT1G6Ccm6hkGeSOdsn40Jm7oCI6xaxE/BIICVvvF6uyooj++Obgn7dxIurNmxctescEgVApH6
azMlV08qJVF8LjJmyltN2MLFgk7zabwp5d7bYPE7/kcVe66Q55Ue4Giw/Vh42Oq55PmLyuwVCrfv
q12Qg/LahnhLSpMVZaipJoJXUyxtfLYmLfhgi/3iW/b4oLCqOe1eVA71k1wCXBwxXeWmHoRaH0vb
uKWbV9dHx5Pc/cLg22Yud4Yb0rYGCvB07bDFZkGhRpAABoP1DXUlukBC+Ffjv5H5fDZ1th+7C8Ip
Her0j0DgqUfAGuvaO17Bqgn/ftq5Pb8fpum+xSGRwVRbY38zVdFf+xQh+uZs9qS8DYCh4QSPUeaR
I97mDpu6CPsV192FZ2WJ6J+qMdk382k4XqCaW+azok3pJzddHBey4AwFe2jcDV+fns7oyhRSAXTr
GBmrhsldjw4T7Fq1hhkS8VSbuoJa37/MWReoIfKAnJpoy3aVWpiF6/JRC1oXCY7je45uxIWVmhhd
NSHikrOf+tzmqh0xOc3AZ5LsBvBsrIdTijhfd0wBHWf3KPfDu4qE/T+r8jzPMSOLV2yaw8c4UhRS
IBMSIa/WQbjtvBJQSPc2Ht7XXS/qHtsqCn0Eo652bdOcPGmXfCPOrXNBuimeZTACRxx9V3FkS8Ry
P2DLVa8ImhkQOSFk+4uVVitqNK9jiE0HT3yUR5NpVZEdom5C6PoA2+Tm55TnnC+lXQ1AFYbqeYtJ
820YTLuO/xyH8cxXNDyUX7H59HbQ8nPC3/Hmc3hRkvq3RZ+XITQAggu8M0viTjeoQkAQsiROBXUc
aTr1u7M5WZt3xluRFZoJHmkyRNb8J2J6priGPGROKZ+i83OXl1jrFB3niIty8f4sNJ6XmlF29iiv
q6kO2WnAHn/vwpr+wt9ggf3M/lkcf8/xcUVwpLO+3N0AX3jOUSXsyxlTwngTow1tRG2WN9IPKpmr
afyO6hAFR20L86hp5PkCmPQ9+lWmnOmj4x2B4lOQ0PbqgCknS8S/rpKp5o7NHNtt4nmCu11B2vwn
8w6D76OxcPXCeVbDsz6q2W2GwWBzhyF4bqtfCPO6QYsiM/aRU64n3IyBknSbCAZNKAwNNDkn/vC/
sl0USBjP7cU6Tr17UmqGHghR+rVPy1ef0h4hCdsWx6LXjcRkPo1hSJwuTXExKm13KcZne+WUwH1E
dXnz+abwfBw/uQezSNT1pOFZlLqOIUuh7WkaP6UpNRgpQ38eiRgrQoJsFAvGItN0HG0APuI/aeS4
p2SxLsPd89MOmKCIL+dW2UC9YhJBmUWShzrqDF7LmqPP2OHkVd7bUBExSm+ZL3oUQIAwo7dqesTV
S0RTL2bCpYtTgY1JNmUZIG4wT8J63hgNEeUyjv284PrL1qPfiZ1Sgi+ongf5MmjP5nqEdlMYZZ/l
hw1l/dSisFtwgyc/BgmZE82y3NqoFXTbavSlsysxyvl6qdC8m1//gxE28Q7yC2PQbxwqGTjHSJlH
PORqfm0mWCaeqiaRUA5pLW0q8M/X9CxCWU528djK77wypGpYnNix9fGn0+rAdP7NLX+goIH068FY
I1/Gp9U1NJABkk4WVCNm8rnvHTjrs/XBReoZYtwLpO7BvRDL2sO/uy1CAy2wUDA+0lmv3r8PMleC
GfkvxdO153Hp6pOs4iLebQcKtUkjaUFAFDoW5Z3kc23oAexTGD4/pWkN4tvAQF0Kw1OJRNaIRC1K
szUoEOLqq9NGzCr1Hluev1LykJ/vU/5xE7SOPXY5pcbKjkfdwhlzvf1xGhFQvt55EA85WCK8MUSb
aEUNRixtmhW/UQWW6YcTsny3dXsMfovkqYtEyWVPo/trnoVpYEi+4eF6itW0Dvr1U8s79ZfdYyrQ
sNoD8Ixp62HpMAdjvnvxFzAJ8zuT6jZwcBNfdDRDtGSBWnRE0AdmylYvpTPU0TD4l3+g1D6MFph0
8JqmWfvEX8XuOJ9JElOf+OkaaNv0cXO7gjCVRzqXszr8H4FszZ6nW+Y9VEBvkz7ekcELOofd0xFD
Im3PhA+KIp9K0ONsHfOtpGMiBSbuciocxsBlKy57Wd0VIikQ8/LrmjLugdjTMz6S6VdK2MVeTaHp
y5+fyQeqIp5dTxpgrAGvPiwy/yscm5W3D00GLo/GB7Iq5LiL0a/A26GdaTSQzZWPuAATw9Yqz2oo
1jITd3fBaMeCepd773jewMXqjY/QtB0mkKy/QbMxkqnQXwkgKDL54VAqR+R3RuOn93cPrneHphnI
ELQqOhidrLGesl8ESXM8PanzovwBiFNB5gSQsOHik7TGkZbzTuipwhzBO78IiV88z6J4RlVA7l+s
jAloZ+oevef5sOFOfZCyJV6vfK7FED3rP/sUWLZgVefkTBMsPGTMM4RCoNSgp3HLcOw4RLVPzq7h
9Zxm2BFFP5No70lbHTHLwHQQkO8w4LAAmQNoCwG9Lq1LXBh3xAWjH8bon/92u7zpRAp1x1YEE82A
PeQyInn08YpiobSWeLJRvAhmL+XoYSTTfNEsq9y+9of7dulk33g1MUA2yUy+TeDwBgA+mRpjcGCK
POxuSLnIugBfYQHp8v+o0cClHWg2dMM3IenICuJ7Xcbo6fHxQHJSWGWJF1Signmu6MgeffyORdK1
kfGvsN2+XQUPKWGFMINAMeu6h6ogsuTvEonwQADz6b8cM5DbBjFCBjMt8oECHrW/5biyefy0UXyd
7ZPDzB9EyfZ7LsG40Bn+EYHZK+MD50ZNqIN63QzW+NnrX7uV0KD4TXuzi8+kos85oIfwXDZgEAGI
5OsHMiFB0G2Azlfq6ZIvv6LyqF8sxrLXVxLum9HJ4xgwIgwHhtF25bRxIAOrk3XZVJzikWAdJ7lf
yY6VYbvYEUxm5ez64sMWHrD+zBwqsr9Z+9y+UVuUnVG1bALmSq6vqAUvY7DtwTP+vueCIC/UGysL
c8Y2K3kD7O7r7oZC1x67zSCH/zEn+BmwsPLRncbUxMIVD/zXKtS4qVLwiu/ZNJtAV4gEp92EpRRJ
/r5va1PjzUpjrKB+20WYoUet5cRvR/83f8ALEZqIFhlH1mDh+gmOrl9q06y1tZaSqNzYRxfJDAOI
cii1K8XxLQq0PfbI2GfYuXkwnsgZbk9N/1Vcgj0q83SoSidGaajlIKdGWCDt3NAU4GRN22kMv/m+
wzU6X8G5CQPoUNjKLUuM2Z8aVGDjZI5+PeDS/WbExaetMIZb2G3RWmL07NkpLA8HZLC55UJJMly/
D+32r5gRQQ6tgsgsXRYBUbo+pvva3JERs1fKsbxsd6a1TnQJ1Q+naNS0qsx38thNMGwK8pimzZ/x
Y2voQk8ktO4uIiUVt6LRaEMVNb8Moy8yq1b/r99byKp8lHSxtmRzvX/uqTCuoU4QoidRztUYS9Ay
9U7xWp6ZU4fUEmiwAw+ccax6kwKgg2SKHKIQNDpGsFlw8QkQpAqUurGpz/4kjVgk6SbSqmA7gVXK
FbNv2ucjg3ymxofN3UERTZ6fe7A+0WH5E2eL9efZhqArbUnHTS8x7V0M1GtRtiVNmIZdwDUSKBbx
t+pKgrWxjnt7QIJIvMX0LblD6nQCYjLooXV/y0GLLvF+Q/+078QbuUeN6oeduFvZ6X7Yec1xZeOO
+zhAkaC+wO/0CFy2Tk8qzd8mDRI74/J37y/r6DFWmlY68KehDnpmHIq6ootX+fFjICI//BKQBDb/
f5V1m6WclofIzY7V/j5P/JheDjxy1e/czFJAhERSnAZ7lnFN4DvvtDsJyGfMlgsz0BYXxSOVgL3b
kQTHUkw4iqtEFpqJRaK4inEqERUYzU0V+qsqJh1yh9bsNkoFww4DYgoqI3jC24IjhP3Iquc5VbzI
W1G3F87P+iobwglx91SHlAm9G3mt/YeEfjcgAsLpoolsxF32m8hgHr2HVv8VepEzZJogoxwjOnBs
Eeaytl6lrfr/iBj65KZT0NngNmriuZ/gN7m1Hgzd3Q7+GfSUWx0kzmGkEM5Sze73Gy+2jBGt3VKk
Kf2tkp6h7bwwWj3NYROFNDbuBP4cIJNDZ+sDS5J3uGb+Zm04yRbNPOD3tm6GSk5bjepM9AnyNE+g
E5iVK7zrM1xGrws1AG44uev39xA5TgxQmBhMkDNOsLgLBXUuUJIk6kdWvzssnGUduTX4C+wtuwu/
UkvH9hJdfLavlb+p9y6FOuKaBtd6ajSg9x677aWIE8JX/+MCKFeSO+XhMd0H8S9bVgTalexRtxUX
E9r/vPDdjUjuS13SaTlG/QxqoPF8bFNWBJWbXpQfDiaGAfhl3VaQ0KByGh7okiebtoYPlqEyX0nV
7jyhPDysODP3BEEbblEFGU3rodo/UayJK3+sSH7I0FW7S4n/rlBu28XgOE+qv9VQwX+R/00GX1E2
C1nyg6H+GYqNVqN2Dij5HIsDvyjTy4olZ4M6vBCUkdVtvgMC49EidLvZZKUf/41GoOF4r9H79Isr
ej2Enwj+o7J0jhPBreF85tYmg5BkgxfrDyGOSkAP+SBDNnVqOg+ysxDqrMl/m0lodUNRxrNgufQ0
S8r1FYSjjFrYIiYQBEm+ut7WpFD4H1fzFFRAo4NcRH0RylYh5Q+H+HZTKQtt4l0cpsf4h6PyJ7Ac
jyJ6Mx3k+MzuQFMFmh4/s+3+h0+bdDlFDHMgFpmJEbQdqjoe7ldND1tADh3q2yYmysmUoHV8A1Aa
t7TgcbVcQPgVE/roUTpZDV+2YO33UHwWTS6tgtg/Rosi4y3qkuFuzUGi2k2baUK6bAQLji6SPeEO
O6komZWCSqU0LUxb5I/i8AaCgun8E2MLPDddHPfYkUaTggNx/VI9mvG574fN1b6UA88kX5Pa1vY/
IwTVOphX/7AS6KUILPcdHIIW6nqOgasZ1tEvaDO2oVO+g1+YwgZZm5B0XAE6bNteadkA0aSdnf/3
+Ao6ER8ySipGCEW2Y1j77L4jqwykjSS75X7c116ZRSdXlPI6Z7MrM3BI1f+B2GgKmg3m36vBGk4f
t8XjWUx/zzjMWUI8EfS8cKgzWhnixovd2xzz4wRMDYfZCsG66O2OUdyh/O4v+y6zSBqdJVV4oPDq
xZvNBFDHO3h6BHWH6j+fsyQj/ExeFDq/s8tNBgFNBdCNuk33Gxo3XIyU0jHYqWteuM4xCQB545kt
KbNO2ByZtP66TdeZfFfYbK0dX0BvOEHr/5AjXWK1UU/j/wpdPIWFgIDBMFDoBorzavwPzJsHuW9z
xcEu4V61BGliEUlwfSi6WaOJeFtRP9GVUVLrJdJcXh+o+a3CjfKh5+68d+aqHgJyvB2KUnLMBBih
NYlBbLNabPaV9YCU5TdK5s63QjLHq8yP8iTqoTszO8qzEs4JcJqz29qJMRhYRSJ/1udFnnVLDFnm
nPmKfff0PSKWptpAc1N7Zgum2tspfu+UAdZh+B1/MnWsJBxBgWn4jB3vTBEFZUJfucCs9hLf3We3
9dTjVygnB5a7wsZAQX3ep0UREAQUKe6FqBL0+gmOW4FxSfNnqELmQvvv8i3Uu0nVfvLgcw9E1AXU
OYrbUqxksx3lw1gw0SBpJJHTS2ZAPMXiIpba914O+IMcQUCDN8vGmjEgNtc2u3yej25sGyWmvV0C
qzLbsqroAhPysB3Qew1jUwCsDK5CyaT2TVVeilhF8KBWth0ZNS3eh3OVlrZStv5MBUAJLubQ6V9j
1FfGby6n+tHgM4nZWDaFCDJG+oSDehAA2aW2HR9pCkXjaZBV/QSKGtlfIzJrHO/YC0WYyQ0m9QeI
H/PBxfjHNSx8ezNgyD7adn6nNEdRaD7fgdPLoNVmOEL47EBNRoRzuohbvH//tOuVax8AAQbJQjGQ
Ra1knQ40P0mWxuZNIB54X62vyKaM+VubSj+MBfx6kyH3L7FDftu3X3Rf9ULw0A29KHVrv6cBjkvP
yXxxqEGI3pLhRmaLVnE1mSIlxKbpBJdkTtrDygbKnAElXfz1BEBfPT+E8ErRvz3AZTPvMeKWCUma
UV3eXj8o/ELoU84VZX5OV0mNLFza/BgvUFOSER0IuuVCbmrxf2n3dGCrxqXSGDhLNbNvZTTuu17a
/EVnkrZ0RpoP+IyPUlR6I/VQ2ukANPpeWc1aDYaFAVU/46a8rIutKKieaUAHFLdkbX1lcUhbjiJR
oyhwGn23QADXYI+0xTkqYi6kKVza/POHRd3OCPFhybTrKkaZvGNNIp1bpRCMl5EBouwRUJF/rBYG
pMHKJHNzURXG7LvAHdrRoVfeh0Dn+YOAvn/U8e5Zw+5jBZuoSMESxPyeKdMCRNG3IpAUfR4ku86w
p7j2WABMi7tber2/8WnRHwSin3fwZygn1DmZRdp1VIINGNGUj6VNznTPJpq4wQ4v/cVGoeHDc0Gx
gbRfGcsNJa/xoWIIREekc9yEFF1D0Nw8xZ9KF14HZzTmuzcKwaYBZneop6Odr7e3qOUeZXm6Mjaq
m4kDjFbQAfmvmh7l32C0C2e4GfBA/C+lNc8wCYfT3IRBeD/Zai5zFsCI4PfVWBz83JbwUm+L3ycX
5jKwUvf1KD5dl14RgyGHPGHGErF/K2rrW8SlFGa3OfTIhL3dRqGnCNkoEmoJXkVKM0o/jAw8/ZWM
rbuITPLEWxNaZ+M5XgW+rCuAXDpzp9MkRgQmMPBLFbWjFWtVEnDUTcTISUfPPrP22QJ8KpHJVZai
YZ+PEN6XidDmbR9QUJLZLokoMV8D4urkNX2XQ/D/qgZ5y7s8zuZXvdUBQG6pJpxGGeW/Mu/WUK42
nJx8fjE1yG9UBjAJVfUmloNyqVwoMUMVeOceHNHUjARgn37g3zSwNtUEk/qB71mPLKbVwu6zPPuO
4LNgoztytWoswOfrRZglLr2qumGWXdNoc9tQQ7C5JhiGswnptuunx2j2owDbkcJa5V6tHdyH/+Rr
sx5QvYR6v1I4GKaIUoJnsBbnWpuVP/F91l6kBpp6rrWGspYuXcTqn4wRRtd3vBWRA467t2/Lb2XM
a9mr2yTa4kEP/LW9Zj/e4mZiqsZ/TGPAoxAJOxfgRxj7Bs4pgUMN/R5pK2khgF2L55scE4mfK7+p
rbth/39xtEEaCOJCD+y3ZYgU1KUwSI6sO01ImyblaXSOD1PKHcCvH6kRoE9kQF8iNfl+opNQqHrG
uETnxnK4rimaLT/0bDnAIHzvhyExUO9KLQRnCq+2JFbKc2eHOb0Bi41x8GoFKEhcr3w+QnCLk2QS
fHv9cS6O6/xYdDEP8D3Oyg5+pM2LyxQBdFQbbmrjCTrDuK89rZ/lr93Mlc7dmFESn0RHC+yHWA7o
GJBBP+l65IUGtIeNk/KfsmZ5FVme6S0vPGrSKerRafwiC4IK93xuedmK24FdOmfw6sEkwjb9YNLZ
Bdg7BR4Mp4BIU0QpE5Ot/y/IAljkO541DwJT5XHsFzRiBIy4hSvO390VUfwLrN9cUmo2Xc30aLlj
TFL9ibub0dYBY23Syn9sUnYZCbme9k8FSGEt+TEDrwSKvtRrj/OPhzfSv8lOugn9G05uudmox+2y
aOSrcIyRaUkPNWEAku8Lf15LNDMKvSqQHUyIVdGKy24kssmEDqwBga5ftMy+tn3GNJXoQ3OJ8g35
Nvs+wkXVWQqHZcMZ15b4kr1ldJzx/ArOvlwuaiuNZ/jil74aZUpS0rEpC8FChN0gcbexWVbPDukK
EevvCAN3qltiBK0dI6dGXfAAP2k+eWeSS4bSAF4X2ZxwYKrrpm/HuAf6HGxCD8Syearg0v+7X0Pe
0tRAVzeL+fSsGRpQ0GuUrwXrbVdwuvb/7qu0DvPDTMDOQVlKEWeXk1vSb6t4L8e6uT1fOnKR5wQ6
szqwr39ZeyqnVxuyiSPbEe0RLLuVUvLSLO/YX+rzEEk/OVFDX6Vo3suzUIgUMHj5NtrZQJHIS2HU
KwVVb5ZE3gsKS1buc8Y3qMQKtHhefDEwK5dSKJL+X1ceiiyy/P0QuwXdzjVPNnW0MJpkO1ynFbE+
5b3zGT7yZf229GclRqubggaukQPtzeipmmRDWb1kozNO9UbwjnSzjctEXN83GF8afaXnIAxDrLhW
AJu6+Bn6dYA4jFDNczbjS7dApxzJmqwZY3Br9QTp50fUXpM+tLLruOKMofSGE5g3cgKZ/v2pBrU9
VAJW90QKF2x/E0LxEFS+7X6l1Pj78hod2/rfbQgDXZLzaUr3v4LPWsCeOsUflmbGGzhtzpXP6/M/
Y/5plapsJzlfhyF12Efqo1VFE1eQks7oK8tdlPkz7+aIRHBQtHb0umvlRzXwx4bH80tXnaxcwBfA
1BhnHCKONi08ygF426HH6GIR9zRjVMsU6itJB63W7um18CRlpeiLF+RWYiOSjpTSZ/N7SN7ZNOW8
E0ZYXWIAKauWk+uuG+/Zdh8z0cgsZs5xUY/D2QuLCcvH5hqIqxeRRezhh5YQ7A/77OpVnF4sTkle
cFXoO1W7PrCMWSvV76PKuPYRlHX6T0km8CIBm8RbDfkBRslTV+KPSjrdFBpnyv1BeEuXx0tkADOX
gG/B7lUAfnNLyJBRWDX+9Cu9VFQMNUNrgdwPv5ihhchL0MKHPqEur8OgS5zlFbQ6SEV6L80v8yAV
Od/vIPMzNR0SVD5TnBML8Wh9t/gqRsKzM+AU/uU9l8AXh30U+3vneW0yp0ccHe1wjvU69cFJvNxb
dEK51ZZUwy+l2lTsyj6n4ku+aadac6RT4C0PM6RC+fTis3u4/Vkx0+HLlpuxtiH5PZq34k9w79By
7yMHE8QPaNlNZkG8aA2+qNAhboityNKgEgcPfqafT+c2eO3169KnG1razkWVLPDX9099X4w04XgK
syLW7b+rqFlCmCJtRALB1m9sph8GufpU6Ry3NUl32AHlgVb7CNDCdvWXAUkHysdL3e7dkMLahuiI
4fX4XLyNEktIjAtplVfONMoWCtfBqTACh5B19UmvfCJLwTCcTSEDrkLAZqwQ+31USN4k//ESPvhn
RNNvy6uPCk6xRFq2SvsIc4sRp9UTkMWUiq+QKDpgMQdOIol3h1N+1qb7AFvaLluLrtw3esmCFHW4
mjwtWeD+O5qSDpQElWbSh7o+pe5YVUf8bXVtZ3N93BFsd5yXTGF/hxZ6s+zobDaq34TMm/jV2ybO
dUkCHtLsQxL8VpK1z2V3cYfQi5fzSOHEzBTtFu4+CqNnJp2sBSoWPFedo1Ui1WwR1UsYUIq24cxL
zbT6C2Y79emr23/HWSabUdWLZhGS3VcY3OMpP4dYlFT7f2GsfqeIIajcWrw7hRpQTwUuByIWur1n
0O7Rv87Yriu9yqg1mVC3cVJ5tEaJxJ5F6tVWCl6cFOvx1NltwGPSCwt2OYVAIRqBpisDc3/eYwhM
Q3T6rd/eSOo0/aDdp0Qqp7bQnZaZQ+2e7HXEbxyTGpKOZVNQPF0E73S1A/+x4hQeEnmvCLMN9RHP
rrI85JEApCxjRr1+6mE9WdFAXfL+DMyEngw8chiyqRnrYLstZC5MhS+lkkk7fcFhUUrjLCmLQGde
Amlv4E0O3boamJYQ+UZHJTcBG9seKTxosdhGKOVaSq05ieG6PzQxqGp0t+K5J0oIHBTavL4dXeek
rqH/GbQCg/pctK/QHXj2M95QdsswgWQ5g9xhW4WkErn/gI0tiB8Uz1fa661+E5flKFP7nR5SWgWE
3e34MTJm/2i0QbjNEROhxFtsgPlEPWHTyMEtTqJBzlHPifKPuq1lqTbL0SgJ0jJ+1m0+zyWIoPiE
W6DQ0Dy3XB6vgsJ7hSqBv4kYYOYVIcuGNbiuZPHZhPw2E1IKeE7zFohf4HRqkdeqB/dUsN6+JLUk
kFru7APbzXlSpkzohubvtuczyiA1l6LOOl7KAlhWLgQYhrLFaE+xWSyb30bO+jst9ffs6yPJdrdb
hQxDRFxyYkReyywl/gQMW8KEqYop16JubyCzYQs5Sbej2ej9Qx6ROH7RiMTlfBouw3/NwOgdD48D
UkBKfxCt8a/ow2lQNhlIkgt8SEYibVDk5o9sO7MDg0AW+1SD+F/SWx04hHt4jNBmgxcBq8ZP9oah
z63Zw/LkC2BdWopjj9wWO9weJYI8LNVcUt+MMWpVDX13lYlk7/4RmCn7B80Z2dOyCmN/f/xw4+XG
lLko5xrO1NHSQnDFRFxutple/IQqYifshE5OvtcO6VTe9KQC1ICZEdyeaPtHMzvqjnsAJcnaZBQO
Hw+CQlVehpCZxerQlhiL1r3T3wKM4b2ha9tZAMvDb+1bXGlpQCmd+xHKzRyb8WIgS/S6f7DrWqIo
8CbbLnXu61bNF1rjIDlRpgFgj01btsup4FnA/2aXNJvbqXv4LWKMquoTcEKiFycaKE3VlSzYsL89
9aR0hlLUVrKX7nOaVEw0FR4vg5U7xO6PfAei9AYH73r/5a+09O9Ur6ejGg06S2uy6z6LhmtlY7dI
1lpViGrHeTx4t1D6oviYYHpIQ4PztcwonryOjowUFRckd/+aWdEVfcJLnTZNl7F+ticfyx6qowUW
XsQlEkcsCgssiMbtw+KeG9Q1PZSdLM2uq5H7y3ktJxggiBkbhWXEN7ntpYtcoamizfFuGIWDDgJJ
1PMbKb1T0p0NC9zzq2li0VVPdiwx1C2QyhBj8dgs7sRweMYWViPvq8lv0QCJcljK+VOFwalZafhT
L4DGU3wzC6LrQlBsMss4RdWuamH1kvAump/n7GI5/xPZiXuTvWUYV8DA3veBKwiqDniYClaNwnRB
a4skV3zh/8kAuum67cOHKi85n0bxcOMN+2uB3DXt4YK03keRQnRZs/Jqk+ebPVmaSjB4gyof6eC1
97NR6lUAG5TYZ3GbROO866UqIwS5lGr5LAlml9InIDxZna4ZTE/Flhv1wk8sytDwkaZvF5qTD/M/
FAliWOs0GncCe3RyITjejWMjfzSgjAt32F7/aSqOqbdlkGYpk+o0C9H6qWqhRWsRy/f0Xk9ulWgn
nRlacMaOWlnZTrVSoHpz23Sx4rw6BWqvooQpANm04juktghjBZ4udyr8AUn9ySiS61JrOUCO1o3C
SmXLimfE3K/zrhUkgcX9mr9/143y9gEHRUTxWvyiWR1xtkvwTAP793wQb/yh4yccG3RgRKXdvotS
C9KS3X6NiRqZtVeQBvBqO+Z8lbTSizN6n/NZITsAfIY/CcGTDoDtcORbYwQtT1/Fw0lZXRnFEwwy
/mfWTw58MbzOdZuqCfIEUFxLwARQ5E6GhruzgoeXRn2GcLxV8tCoo7S+zy8XXosxmklIRuivENMy
0V+ruicyMblsFptSX2rctXnhuck0hfq8UAQRvqvZ9TA7I3Jx2DDRivsLPN4bdqgdfiPYrfuv3Bfe
tC2+4SIP9SXgfTGkB381G9GDMNkO3f8YsWEDtu9iPg9HAAxgJ7Mrc8PEc4D6sRkeiITGySQAI/bU
MHzjXJ6T6s8bt3LrTnl/jinr4AKfT9sPXzgvJSUl+tgxQijEeEOX+1I0KmvVcpBzcr0KkxkIb0n3
ojf4lri3PAqwlmSm5E6tW71S4PH4UhsfOkBN+tOUvkOyHrdHumInawprnYbTi9GiU/BLmTGFjL8w
2Iq5MQ+xgq3JHMlQCjQ2T4kcS0x3/6oWzr+aVHKQ6i6hMDaGj08gS1zfegYo7xySQQLaHaadD/Ix
FloDUTsQZ5enwdbJpQ/E6PKxPe6FZaridRS6N8SFJQVfzJp4r/2dOQyV/ZFTzKuEWkwocWHl0tNr
HYhp4+VBC0s2uL9G4A7y38gN9hDZEA/32Tpg7E2ZpWExJxWsMwZ9HbUZL+ouCe+TAUOcVNunQJuJ
yq/jeT96rZCCSRt5sQvfsubiCy6ZzjYTKUViV0UP42knHKIq7oRDFtCTs11DqTVKTmYA2YI/Qrj9
MqJMdoC/+3eBDi6ryx6VcyUmbYW1qSysS6jzMazW2HwchKX5F21VKl2EcOWUw6A0CFrATg4TPj1f
fmaACUcOQKsPxiGM0Iy2HW0o4UTUoiw+/LIEYUNLGqhIFr2AoXpzHoF4Xqh62sJGOnr+oZGtsj8A
0OuTYBl2BlwwIAjUmixEHnpBtiGw/nxAR5ZqeVxWOufGRPoc9nqoL82Zq9GROSd8HgSqpOZWz+w8
T53+Hv4R5QUDDUGZpCrT00ATs60Wh9ssOTYmMYOk4Zoqau4vK526jHfNWvMlEMdFolHsHAGNmSj2
+DQS804Hy31S7fMceTbhAiUHy+5MI4tpARH53fkOaDC1a5otvJDz+segUTa97WnwhestJ0sdHdHT
I1kxm9tfoLe6alYZRYuaLGymGKknP3r8pLGJ4FNsGdPZdSze+PgyVo0dcnv0wTnLZ18QBW+gFd9A
UwwMyqcAXiSKLiauSuI/tlWaOsj8hpSOrg6XE6/JRBWr0CxT2pF2lguL8dMrzYhTwhDTjhKV0JKY
mbFuB2RG8KMHEMioNQCpO9wHgVNQN6+bQnIaspfe9LlmAEVcL0+M9W/k83o0iyQ9/mLpnEjC3uD1
NMO4weqbjqmVUC1vVQKzmKQQzsZ7rUCtyuqhtCPPPcvbnnsRHxi14WspMbx1ESUoHJ0JjwBTrBBw
uopyLSOUgwON0sP1Avxwo+Fx7LUuUFbGIcIVvPo9GVRhiSkExOL87ilIQFTXEJb/01ujqxGvNnxA
vO7tF8FOTSgg45FP+3FzhF7YO0T3e3oNtyl7xu4kCcWVrRU+rkd+3A7hU+3NaD8BULi/TgnDniDO
ZqETpGf2oN+e/QZSSM9mVJIZgJdPCSuFBPIJZzWHjmJhmHQ/cf9lIXZXonL+0tH+kYKqAJpR3WwR
ZFsdYFJm8YQgZiWk/TtzTcoUT8nHjA6bynRvhhbl2tLDZGSUkUlNLeXyV+14SidbhnE3CPbUqt3t
Gj24nhRA+bwGXOT1LPxtyOF5nXHYpk+hMZYyDzamw4u3wgVkNOYd0yCsJeIIK1gwxkPZdiMC8uTH
yJpK4+WZcCHvb0PR6P3q5J4bAceqGZbulmx4VGKXpD3yrWwih9vEEdwoiTCbigiMNDUp2jgQDocw
UNzHTvPquUWKcvDr0M8TXPaKpqaGoNYMPP9l+36sflO1EKyNAANs/ep9ytW8F+lhnZ9nClirdKEJ
S18RukPjcuKaCFJXzTpxCFjxkaRP6idhsKxGmDWWH2sej1SbKhacArOnH9dJ6c+n+ZQmQed9Pcr4
1SKY1J4tWaewx8cReVE51PEItNoB79gMNndYmNMUJRPZHI58G0PmUiIkX2CmK0wFeIYtSOMiBPZb
dQPR7SLOEVOgrVgyhrMpC/sCEuVTV2bGxeduJrOzhEqGY2LFt0i7mIbefHLlCFA6lZ/N4g2XILJT
/XX8hxUf7V0U1L+G407gYHdpZ9PiBGlwRahMpsL6viEjUYdK0QzKfe/k/zvywRX/vnS2DdT1KTWn
uGO+0/qWQTLjOwbmz8AhDxcjH5uR5Xu02ssqoyXZVR4uh3GxSuCMjV4t8mW6qcNRWghIjNg7QZKR
8QoX2EsPOUHyUiWQWqO84lpxoKyayMWM6WMm6K46RDMXqOe98QB4zsrb0/FvZRgfaTYiV5CH4gvq
Iu8y0xQov+KmPnGprRakcMPEu663B6RqJ1eWc4W4qu5EIaseFy4cr/MaLT4rKC0OQktL5cIfs7dy
ytE6F04sUH0S1kkYmFQvlHfVgi90NJobwHeY9cBSoMA8zg4rtDGIFs3g8u9UPVwwySZnEQq0olyj
zzmDIEes0CeRH/0mL9P3HkIrfxL8oiI9PZ2ooYf+/8QIN+YuyzLBuYsGaYkhgNdUn30GmXjUgCqP
F7QWbPYLn3eVhOOgx/k3XdziUjw2FhhzvUuHBPb5vf1+JGWl2nURj3diMoMLuhUP45alwuJ4Sl+4
0AWZ2DT0Mju5NJKSf1yhUC9Irjd9Wv+TWXcxk1RNjpThOAMvdZqHUc9a2QYblUVJZRGUF8heznvT
V+ntFN56TjC59adGIRUtpwxzCJSG1VUl+oHbWqmF2QSPcDl/mB1r0C9ozaUwppXhAHKqIekt3l67
ivtRtv8MwZDIkDzUgBYQdnz4O6PI3H+w6ZI1qyV90ZN/seCeu9uKz7sfaamyMBJomghvxs6EWuF8
1GrMNf2Bkz9xLaaSZ2eCjm0Wi1xr/LPPuER1I6eLPZwo8LBILhKLRlobUEb7uMS6wMdk2wgCHArS
FnSxAFkTi66DRDzD9mJ+kWQ71Vc07HWaC4w+q2E3ezKmJmW4G5WTYPCymU/fIKpCoMc7F76lZHTD
3WGIcdN0jRgt7X2EptqV/hA52ktecKUaHWOkdwzA5eDXVpgid7Ew/VU+NeNOzwbWhu1FHZfJSH5K
5/k/VhcJnxr+Mao38urdxOWIpaJEvO3qwfVFmOyxJSLg5QQAJwmvrG3HWne2r/HJtrQOZFpJI3t8
Bd+8ntfQTcgaggyIuFmRLKYmmxK3AejhaF/4gEem/IyGzzeVcqmfmH1JZHiRgQD+I30OSdn4Sx9g
IW1IqN0XA6nR2S99m9r7r1T/caGyEQTJUSiQPoQf5d8hJ4K9waRouG2myFLifj88L35E47swGpAe
jKpaU8539fuNfxNiiQ15+1jXMoHgAtcnlLFo3R/ktoSSbKCIts3H/UgXEZdt/rlgeir+PwPbsGHJ
11UJncUUJgMCG49n7/S54NP+0HVaKyDng1uu+0S61JuRF6hFdWsZfVG2KcE8NbvOklMdI0DPP78F
CBwiF6uyBCI1ilOYL8lMXJceMcKM5JjepV2nxCJoe4o8xfTFdrWPaWGbyARey6sxvd1oAqG7ay+T
SYxRx2yDaQOPOnCMs0M3xO34B7LPboGtgpx9Cg2m91t4S7AC2jrM8YvTxPrylfAd0dtVdzEctKFe
ntfjkYwqtnohR4jkVMZDucZutOQVe8X5to8CApeRMtoe/Lb+nRqn1gzcawBCR+X+b1qMr/jqMcLe
91dtSYA2DlDsZ9gh4r7dQIB0oGnCDHgeL36Xivoyb0X8P4/YRu2rqGU6NxwY4084ATc+jhfeOtvE
tRVdskU7qm9SpZvR8/tWOO8en7yTJWw0+NCsanQc7wTchYZlVR/bf/h9U48SvpO1mlbiXQoSfohC
ea/y09bIodj+Uk6k/wqmh6+NQmpZuW8+74VCZTL1C6Ne3hZNbNZZvrpZl9v5D9C5H/v3lV9Tv2kj
EP5/Ok1O7x24lK382tatFNsp9rXxO35OliLKLxb25BtBH1Hedh7v1wPI0D2BIs6v39eMbKYk7f3c
UTU+L6Wx5+G/3Or3gD+6oOpSFKhKex+iD8CvpNrADK/QuZg6ncPoJSzsjbLv10HYMFs9AINfuvqh
hXkBnkr7BHY2psOzXcuOmFPwqN5qGjma7TUoCPvcmY+q7tvYgevhvSs+S15LBnGWPtjSuAzszO5o
9WLI14yQbnSE/8kwIOIvHqvEyKgkFgfzTiLzoAfi5ztE5NxXE2oOKWf9YD7qAjo+UE1JJ3bLbMkj
l6pRAQyfMoOlB0Bmux5uN7iC9RXXYomX340mrFuEDFOyk2XE48UjI6pGVqvpiZuw0/RwYdBYqhRM
QIvXRsInr7LFnHPKXPYqgjJsBUymjWRpiREwMZS78qtdP/C3/5xSHrU+nmPAy8cSQy1cbtx/RU2d
K01lqKM2FEMdUBahLF49jJCHfWkXC8Io6rwlYz9u6hzTjLqYLIMKCY5RCbJfzHSK3XbAkId8zp2K
jYhbCpCFoXhuThnk0zrG+RlX+iYl9tYKiOV/87Ly3DV9XiQ3s4AAEQFrsghvdIpXdJBHGDx1+hMn
As7rmU8Kydrss7mjeIziqXFRGEE4Ts7/JiFnWcPdwswm0UhCJRJLkGOnTe1RBgz8UhfKgMTi5UjB
+/V25udt3tIxe8ovIORt7KPC7eCeVdJJA73D0R0/dIyzSBmUtmZpsJh8etSEqZFCfV2swXQJzX3l
+8YFGxYbQ6evWrPYRPkeXm59IQKVmLiYQuxK5zmbAp2he1lH1/MVs4VAzV5byyxTXq6D7Y5ESP+Q
n5yis6kJZ4rXbT2/IouNj8buToyEz8DyLjbaxjp/L+E1wIF/krTWQTjOe73Hjv4tGAs+KOVWRa2z
Fxq/hVMVMECBgyWOTnyS6yZ4qhWED0V0flVkPNVWebOrp86k8CLTLXWBxj0srHsE6FvRgd0dKhQ/
yqdlASBauhCqaTPfaiXDE/6AHyijo07SB+nkTItvEfIlxCylKb0lP+DdeFZPscBnYnX7uuT/oWBV
FndXiPULXrQtO8XUmXCRrQzHOIamC3vy29IJfkk/bQWIgQbgS2CHgVh1dR0mA5cnHP5SiPTR3IlZ
YJbkSCnwu1q4B1HfTVuK6NOyzYrcHgSo8t+IQ5IEwcNig+SIjhM6DK1/Tcn6RUvjUcVlg4of6Lsa
/J58UpcKWMk5zlDaQ6hhPD75selg8CnO4P43LWp1dW8PUhzh+wvW89G+eBQKmInZm9PSAPXoGVhc
M3lWYy3h4IpXiqTTunhHff6KdJOMS9w2Lw/zOwuV6DjT290WPXhyXFZi9oRnqCPY0wlSp0c5V5/3
2vtDTb89dJ1V6lmQI1q8vJJxaDQU94vqAqWEYVMS/31o+//icpSCnFwhE/eeeHl9A6ShBYd7038A
a01Z9kJty7UsWsknPmBhp87SfBf/GNsN7SWxo8LwiKP8gvwXCq3CRN+5NMNFABMrN+KWvvy/UQ3M
no/aOyQVrToX+40O1tfV507BEESNS6KeIfobpbtJzvGU3Vg8q5PO9HOcFv9tRMYGtwLlMi/pdXfK
mZ2NUBOjZXPE4bheVPw8YBu6GZu81VHA0vJ7Y0Tzbswn0egVrGG1OpeikjKhgrNQnQjNlv7hpbaq
Y1B11ad7A/ukUN2oMufsKavK2NX3MmxcbIjXmsr8fM5j1hVkrBrdbj680vMwBtBRCcfJDj0nw63c
TYyhee2RDOgjkIEYPURcE1qOmWP0TiBj93tCbiXbhnN1RJ5cseVtmbN/6XoboLINsQlTFu5Fcwti
CPN1r0I2vdfc8P/oOoyIHujC14vI1Bk6Bs0RyQ7ph3yE81xwiz1+s46F+Apk11qBLK+hbV521g0A
FygKF/f1HF8pQj824P3JdKl70uEQge9UfacRGbIAN+ChOczhfm4XN7U0UkFq075vZSzE3PREmTu9
6g8wztbyNcXwCTlKooRNH4eC3q3LH7yIy0/Z2EZUAGIK9ukL6yFwh+zLK5DvGF8ltfGlFaez0fVu
9ihyss+Qrxy/DahAgmxCXL2OYyNAjG7zI0HWQp2TuURTLT9NYM88okCB7cmqGOYIUbPMG3xbkIGA
qOdrUygWTX4432f36A2zr93GsxUEZ28mFgD6xzROUT2w869rKbz08n1oMZqaeI/g3l+GfFbLRyIY
cjBa4iHaqxmMyVczNz39TD63tPdmucHLueh3YDVj7l47vYvv6XgzBfGeqmnw2svvCWddlU86RY0L
qrlamRMQepExmYu5P0tAJf2KqVF5dan7CBQAT6RCLStu5RnWPRZc3uctYcVgkE+A3sPdaXhE2B1D
eV3jNo/jH0Wgy+lEHV2KZMyucrMSiDxnIhmpixWWGFycZ5lXwFa7BTPIV4Qewcgf+Jgp56X3ja75
f7edyC894WAPZJ1cGnpTQzxhcVsEH824nMiSCBGzKhMkCJCS5vzSyU66XyL8CQsRuLY8jHK2Th6B
UjoCHVU5ni2XX9LyRRfwRbhVvpyiLhPv7g7nl/5Oen6xc2Pj2nEzHgChVOBfSzsETLnreolv7jTx
M6Ev5eEw9dut2+vm8ftbQAONaNLs+nnAArIf8YOUArcw0ZQX45NQreQUgCqYK1gt2QZOqRQlkzyD
yH3X9yCsnWJVjhCdGOfJfuFGheKqpci4fTK3bk+Soim9ru9IeGvKFb9OnD3jqZV3tIBYRtZg5Mid
BmQx3Rjqp2UQqfOs0SnBhSufP3in7s8iSXrnYlq1Tb4HoQCcBeQ31EzAiuaNV+O2/+rw6gHsouuJ
Lco1xWbONjlwv/sSle381+TMj8JaxAYXCIgmpJ9yqy7vKFR0q8tkPnKgGizQtSxEVVIoqLQUR1Ko
P56oZhpGCZX/wG52q4q8d3UMGitqUmg44tIgPQEW0vaHODGnJzGGM8WSRWdbKttsqheOZ2WwW+KN
yLB2muCwdbjBKigXwgL4a2o0D/cz033hInRJZ8pKr5sXu0JBU38ZUzDCkL4QnCXQ89MIRLtIFHfp
lWxBx2XOhg1R6M9K+C5hnvL1F0M93B1CbEBmREJ2DlSvvfSMaBVQJaOga+yAGwK4Kl+76ldfBlCP
V0MOqpyJzvBFgqMiadnVJ/tNMlrHHD+3Frpp0BUXr/jcfRtJS5t7d+VsXDdsHQztKBk4wOk0HOlm
L0Rz4FQc3q9aEAW/tnbIJRe0c3fkleYBtkdZfFAJQ2UhCNnELM6WMbwVuJwFK88nxtylyLFT/Mby
wwyxRsRzuvN1PkvXoNQyHIpCQnNr/SFVQrzcU0jxbziT5bL34xLg1RaYlNNFxMAGhXxuZ7vyMSeN
pms2YWG6DCPGqMiKv7z1YNL7igjOcgrI80vIIsuNLYVx/lSfEa+uj52jOJB9khNItFyLq/lX4ih/
rXCe+rxt5kvMgmjSPbCp7WTLum9SMj0E7s08cinfoimB0iMqvyx6W6VqGzixadPqE/lOt2MUlpN6
cvz3s4LBgv16tRXZc2VngqztQLgJJ1KrgU507goC5r+5Y1rOUnkk3YrBccYgmzVOtz7Y+OQEL1Cd
WZ3ZPrkaz19wxZAPRXmlPRFX6mjZAiO++3HH7H8j7eB1MDgQ9T/IHZcn2Du/K1nfJeYu9SfTN1S4
fbNWjI6h4sXYB1TNjig1Y1Aa9HVhDwkNUAEn7knh/PgJxeI4iqTyxZasY69x6SqfIZTsiL7JAtGc
Z2COEFegHca96VZRGejGbRSgWfW9vEzI/ft2BpwMVf8D2LfmjKrL/LFWAJPNfDko5LR28U/aBl+J
WcxcnzCykB4UrL5SYm0zZCbsHrTDhcm9DqP4u9bF9umPROWDYvMxc+pBS6KEgvuUzGoG/l0/db8K
gpJtewJQLXLXuTMLFvpS0cWZ/LGtBTIumfVEWmEMXEvbNXd9B8qZmCHeuXjzjduianlqfxS49nSH
BP2mYf7Bf03ZF6013NmoPXVJUZO2lQiaMoIYQy/swBN1S9bJGcjdaeleajEjdEQ21HbAR/JsdVLJ
0OOYkAcFNrfkfleYf0smCbXPRkL+2K71VSb1k015b992HuAveaCKZ9ysVbC+TaPu/VrILMRItrZo
rHfxraraX9NDxg6kdKRjQqrtY1DWqXz/06fpRAl8OXn7fV065TvgiipdQHSs+1/ka1OhqNtrU48F
9UMhQmsrG1YnLzbO+L4APUAFGlQJjnS8Lhu8CRHucl7hNuRsCPZGy7lGW/xtLX65fHy6j0dQsG6U
YMwteoQHrQdCM2RaetLH6gcPhlObO8x7xZUHBLQsLPKK+gd7nGO4Bc3MsM7C2Me8Zr26yZkG0Lrx
1yhZC7hwRDr2V12Cjm3yfqQjMXR6WxAGm5qum+CbF8pYhrijq982Kns144iT4By6mkpjeeIamb6N
APpAfub4Iq4cu6H10T/OLrvMvmk0YgYUTcusSymKaHgs4KHfIh7NMoKlAcOn7ZS8HPAFK8a3JB1H
gokCsQKwgi77VGPfEEEXm8DlOWCr1L8XDd7TnKu7WVlskwrFu8mDbqpTjX/2nfSJyr9nvLZcFCuq
JUs7Gch5F8Wmb5tGxSMxZRzmvOZ/QHBUAUWGqE1uJCGzz7Y8A+rTwa7JZU6zE3X84vKQtpdGPIxM
gNxUjHmXqFs3XPx249MAl+ceMx3PZenQsRXEdLWfs1uonlkigM3RE/Z1fGoYHnNkD11ia6+ktbVk
AR042LKAR32sVgG8pvNwtbgATDXk4G4TXonlS3WzHj+ucKo9ZGkaSzqaTSrCw7cEVLwFybX8k4kQ
XrTDVxMFYzA0AkSHidjqsFJ6IJ58uT+BzVU4KTqYtlwFuyA6as9fx1H96hWV80l5Bf0TDmvsx+TM
kDNBUAgEdoJ6AtdnMu+f13h6g/fpMSCkr6WxW4NsXtjclLbZuqQw8Gw5VQ3XtzQfOGIXPhSDE0jD
KWPf3Q+4ib++nM0Pi7x/MbItRlScpa7MVg9n6r3UFfY7imFakZHUmpBFCAeLClKBx7601JtwCDwg
CNAjlYguIc7I7Vj26pzWktBWq31IC61v6+SVkG5CU/+G2OJEYEgqkD7H6EBzuaZV3DPS2ozPrmtG
ch9cFLPrQaH7Kml0oj0RIez/RbAaO5iHina0O9dtRGWVgev5mZDOEGHBdjKWEGkHzqVQMnAKibL2
h/Ge6UC6p6STEBuAf5svgLjLEpt8bqJkP/BHuT6cy+IJSKR+6mvqs6taumi89+R2Oqm620uVbEor
pRIvtPM2bZBX9GTK/1Q/9NDcK8ZiDiY5vQ/0lpIqmrpvq68enLjY0vuvdiS8pEJwuqyjBVY5FMRK
MhOPDWLDi6pzgdpgoGqzxEkh7Tu4nAoNH4iIdaDAvR25PUB63OXNRx7awyEdMhXuxueqL1J+WdqT
yNhQVVvRXFEUrW/I6gJ6sBXvW3eKXJ7+gx7i+w9cIvpczVBIuf6SiQd+AMJiJjUe/UdlCKNRJdqT
gavvC7sNlnNX26EGGe3ZzQBQSw+lvrDjLtF1Fy03aRpdCx5LlAg2ep6P2GOBPL9OyI4r1frjH/gH
7aBxyEuepDFQtEu32o4FZrGtuAAa/l3l7qVLeJaORXJeHgG8PxTMJYOKqDtiwmE8sIhEUB5LCc+t
798t/vpAMn7OrkuG9fil8xnEhf/V1gfJGUWMoKLOBqMB1WYySwAcCghe4Hjnke+7XtGrl5dmNyB3
c/6rH4ukaFHjy5sHMj1VOqPzPwJFNV2unOVMQNbMJhB58UUno643eJQlbCwBZnRR2tF3g8dI7y6N
a5eBHD7m3PN/895GxkVEBiMpomyotD04QICghDTNb05jt+QJcimTd+SuxNt2uyk5S7zMXIb25GEb
UrGnC0hqkM4PUPphTNCYOxg548pTk+yYiqVEKEvStop4+SKQ+AcaiiCPf/U7+UQ+v/wwjO8YzMKy
Fj4XG7aELlwxYfhr54OeHMhr7Fn7OHGXY9XTZMJquNk1fy5QqsBEamRYmecxQpjWIMgEHXOz5Rph
o4V34ektjgCLdC1GsqyL8kq26TBKiWcHcloCy8Chx/lAqyvOHLeMYPnbY1C1A+mwv2pC/S3AFs6L
7F0gE3D3GfmYxeJFqIR3I6vPZ7WQD4Iua6Cje8omhr+zYUHu2+HEuiYtwQ0cpTtPmh8+prz5a946
kZOQ7OgpoENo4t7rs78fl5dpVAKciDH5+ZMla7wlqt/uCRYBTV4BDblsmeEI15V6ti8XE1rjSRFt
IdhiAl+ML6/OOzQOudjXZF4aDV+ZpcunUnb4npkCpZl+plXVcM97Y7vnUwFzWMbLP/veHNFDwWE8
i79/hy9cfCr1JLMDJ4aRwK7DQPKjkzqDj6Y7/sc0CDz6o6sxZUPHZugTTqIewdRqbRJR7vawGopN
AM4eMloG6I+do/rcTL++lKlawzsJ8Xvp53/Jsh+PcY8LUZOrdCrZeOpY2Ohv0H04ZxL4ina67W9m
sMYHD40ZHCOrL6JWukQunKkB/7FkiOwWgENhY2zy3ZKRgvmejm7Ug0Fmj8Zg7U/+QVLKrLA8NtwL
ECYwZxR6WOnJ94+g45DYSDetfu+23xIDsB9Itvt3YqtxiXGxPCXrbOjCxI0K5WtQC3A6dFLd4s7C
o4pGFCahTJjt8k3Kjbmye0yskYcGbYuTDTlsdDfe/sslzW4esnCUxRURsxjKfAWKRkWNNkeRl1Az
+icx9yOLhs3dMRZhWl8RdSav3c2teiDJkILpOzgYcZcHyKXZJD95vYYjmQbcqX5Ytc/+jE80dIOx
valtAQFB9NL2wfCWyP30qVru5rVgf1VUBpY6NcmBTtMGcJjz0Kk6UVBX9RQpwtAL1Npdbvi8s0Gj
rK+dUg7jtF4MGmwyg+dwyqfrvNfAbXUsSWf1tJP9r2GOE6UW9PMmh7mRhYFOI7hWNMbu4hejiRVU
6/RVxsrrp0PGMP+3/V2Nfs8hLaR9wCXK6j6x1JQDJkl4fSTP8P6SnLKHzrL5etsI4Z2rT7R2KvS+
DKGmzHUnGUOwlmbtZbBjyJwrUdOrF0qVz6chaJYZdol8sTqKulzSOMjuVSJLtSD5VWGv9fx7n4np
r85Ru8u1JugpeQ8rLKxkIaYSH/RybPIWdWkHQknwr2P2jZQA3Q0CrMNYSImlWUmXZI+6dpkzXCkU
W4pm5i1niPcX89JQ1VYd0BLM+C5RD6xv+ZkSQk+4saAxiry3nVoH4y17Hytok0ehAIXQpjwIiYHl
rpCWXUN70OuUteJ1DjoQEWkV48SE2FiFuDQf4rbGI1zRNuCHG7hTNM7Z5tutHvWXOfYEgOTmQ1qb
CkKGYoxdyJ9cCe3QkbZOrXTYGopsEdjEqO6iMw7wVN1rDA0EQR8s9cpkU4YN6U2c+5Y9MyQlTi7X
7S89T4NkXKsFA3Jx/mDanw5aLDpFjnS2OWBmD5pVICdtR4N9jLEHSU8b5mYVQc7XGgAeJbVfi7Bk
AFYRBcYDiLIeW3R/5Aw7WpzN7ak82EE8uZPstI0sey7RaB7WjX4Aq6D60Yqaeue8W+A0RRR470j4
usft1Ar9tvrYRjscqnm6O2G94tL9DbQAxLAWrmIinhZskcMGk8ZGzzSG+io/9Eb8lR21VnBYJue2
kM9OwCAUqEKz2AnhJqx9D8Biz5tf2ZiN3Ahk2aqVvWKAlnliuq8mISQbxsY6nSl5ld6SZb4jsp7c
iKw07grYqfKBUiKHojKj6Fk0DyYsP+shfBi/BIcfyjvW3gMS5WwX8yohYDtvPV+1nI6bJ4lP3stI
FV6HC6kSXdREB3QVAxIubTss0ROR97+gi8XlJosqb+lES4wwJZ3eNO8qg9ZWvbE2Y0GJvN91LznK
uPcdZUmBkBrwCUf3wMxyMaEeOvxKY5siY4ydqBaOT54B3szUl34SmiEYVK85Oiq3bAAGMCiQe5nT
guZrvZw12ubSKGmyjnhhYQRnQ3i0OfUZ0Jcb/2mEZXdurdFCM+9MoQAZX0fwh/rM7IR5fe8gsYZP
9Sn91ElHuNUdF365km6u6FsIdDPcyQqVyYkpcww7EpK1mCJBflvAb818PxKmGsaJtjIMmCL789JF
T7tZsnjy1tlPtUTmbklnQpoBCsK5Zy2eqr0OablnH85c7XIWDxxZ1zt28DM0oRpWjEer9BSw+PqV
L9KQrSo77TNDzdH0sg4SONH9ePuayuoNrvCYM2hwgf265dM3ijlmIxDEayVhQTKGqSrBV7buSCrb
cH1diMh4deWc8C2f6a76lUsVVDBWLQqAe3CX54fhw+sJu1vCW9dzn6xkA2Z/aFNq+vM0Gd3xQQ3K
wEylb8lPJ1rP1D7zq4mCGyfsXKMpOcZp2CU6zIPyJtL1s9abZwBhiptZtcHm/kv8jzEZqEzK8d+a
ar1eFzNBJUhFpCrZ8Ap79qJqr09oXGlz+YdPaYfHZiXfK3mYUcwS02Hc7FytPCvZ9u4ISH8wL7Bt
3TEZ0nP2ZVcP5Cf322gRpD1xpgLU0Gm0lLD+IFmj3Ys3LAl9VS3Zaq/cJqH5Nu02Ue1jylHzrD8o
3Vqq0tSTt/LbjPQunRmJgy+fp+G7GTHeFAE/n31LJ0Bm6HytBEgGE8O/lgctWlOI/oc7FHMQxLFU
ymKM8XLPg71+M0C9Vwx8bEIJKJr88Q3iHNE0Ly/GgcvRHt28Jp80skgxBmd+wH54HN6PnC66MyHW
TeIxxOzvWwswjl4XtlqbYA2s6aK5u1T0ZanujfznAD7SPtFCWX0NjzI9q9Dkie41o4BD3elJErXw
6jhzg1m96K6GkYWDTTVuEsTRIoeZhoOm2XO+tdwSWqBYlCxejh+dtk95iI+uEdo6g5ZxutO9sDV8
TDUyYRrwxeHuGHRI4FFvV7TApV7GtZb3uESodf2pw/DL89SuTcG557uRRxYNAIb4AyJ5auR9G/9Z
LmG9TcAMk0qq316apYRozAHK7EmhAFi1jZ7pyqR50TT4Ltjo9wk2MGvYgUQ/LPhn5eDC4GVk3Gk8
HzKSDve7QcxloihG492XaN2GwvumHUSLHQ8vXbdDOlzxQx2/xFSZv1L3ZuzfU2v7ranDeRjebsKY
zue2s27ely/FPjX84ypRi5UkJk5ea6/o6bR9Z2u4gZm/2oUOwk3AIM5g19e2pFp941jjWfflK2ql
gzKxLMpGoCfftjWjcV8G7vTiWFUBw5Rxv12Aof3JUSUP784LMaVWJJLPROggo1J37wWgAZ/4qDcN
X1U3pQ/bftcEV8J6xysjLAgYX4ub8ModggVW1rq5SULcvmb4zb2Zch5oGOd7cHoaqNXBSz8tU0Zk
i9HXecteLNDitZtSN/lXFYru439gWyZvEHmO2Wk2wVg6rrZs0EV9FJzJe40x+AGm/wfo7e+bPwiq
rohguNelCh3RQ+AOusDfAqiFo1hP9AxWc9ETOKLhTmEzvU7qp/fAC7KKUoOEMgQZBH8p/iwYo56g
l7ycIlwS2lu4Z1BF31aklNITf+a28ntLuu9qzRSDbMWGIgrCeO8TFmseQS4wBOwnwX3rz7cz0vMH
1LT5QnqlMGFBRl5HMJIYfhHoo34FeXYB45afWUb173FAhqqNDuGOOKqvsHXhoYkvQKrhPhwr5Aev
q6Fr/AXk96GW30ZN4cm4kOf4RqS95CjNie7kDuCkKFnkad38xio7OcMqX5EaR8uVBw8QTBTungi/
cn7jN8uCywfX5L2tXYnyMVCMblPSDcHt2uLWp/U67ut1iOrwjwA34psDSKaOoA+ShLga9tDyK+1F
jLWFSLRYAx0P/N8VzB79Ht+VSPht5+4dErWdZbMbxl0xfghFjcJUu3N7ExnHu0LDtcHBx3BmfXnO
gV/T8NYbA3eYKtTtj/Q2qT6WNyAJxOXNDxn7xXth1egvbJuUvE7dgrWeaEAjxA6Ulq5UHn7f+1pO
emT3cdcwtqYoF56mg5AsBUEdH1GOy2Sg+Mb7mP4kfMQeicA7c/qp36B51hptr6InIkqO82NjhZg7
niFjkQbfOxuih3hgERJwV5KyafQ1wSnx0sWRDWG3iPOffx8OpPPoQSDuaYmQR5rjxjIGEadkddrf
b1aU+E6w+Ynk3GVgdEMa0e4gWO1ri5K3j60fItFVL2Eiq4T/aIh+vQBkUaLwgHQUvgmL09yJzIkM
o58why3QBLValEGXGmYlRmz90JPCFqlfUP6obnadK35DM+dgxPV+P1TAfsewEa/AlqHuN+WECHk2
vvO5FxgCGCaKak8QZNsyHHouy4PZCkEQtaJOpyhjRfvKu6FIPptqHLF5WdNmY7Iovkp2BccbXuMZ
pYe454dU/QVBZMBXFSE8ebYov7gmY5kzm957MOu7kOa2QxF4Y7SL+AjE68NTyuMZNEMdyjLmG2qI
b86zO99U49D+Mvy2y2H585+W3B1HM4sFpwizCmQ6+5tXbpqSV4KIsAPka/bM6TzZt01mN12H3fDz
svjnE3c/ORp02/KC3zzoV9pLNF6P69o5YGcqllft/y8f0xQIMFSCUFiJQoKjcVxmb24oqZ2NfE7Y
5S+VNskqGY5JZk/rJnuDc2T0VYb+QYOSoyA8aGZ3xt22zScdBpRiZ3dPqXOkyVcMq1CBHsvh57Ya
qvNdm8LRrYpnqMQNZAtolHtZet4oQ83xu9KAm9E2ddrlKnPeSMt2q7QI6m3jFRYvSCUX/1fJcKMB
ByiNbU6t04Ex+FiPtelSb8/2Fq5sQmo0IEwTsmJGAnvDiHuPLEHRnRSMK1jmXdRIC28YrhaWoCX1
+kdJDHhCzZDwtj5lbiD+WXpcqKykqBje/QdTu3NyD+E9rWsI5bGEU42CqZEOLMd50gLPxJiWVXLJ
dx5nrFqyN7TT84M0n4jmQwfDPH2UX3eRdU/D1Ox08m1jjziAmdST2QwzelfX9nc3/oUWdLh1Pal9
sE2QUEk5//da1dWM6VGG9uOxaOpGtllp20VO7+Azg25f9qndOwLvCLigthW7aoxEQ0HBrnDH5rid
TNrIlVv+KXiu6wPkBQACACLu7GFSMPpJI+TjnEHHzzPiElqqlCc4AO4+8kkbGc6d3C8YIskOH7+e
3c2D/22tMvPUr1pYqZumHMW5Rs7xKvh4/YOHodJpyFfcehGA6rVUBtKfRbjM9Q/FdNo96R9ETC33
8mA1l5DldP4xh5dsv9KfFiUrtinshu9hIr/ZQTsYpot/VxzhCxoZ2NrZSa7p3IQzTzHtCuSXiQTx
hONwIbc06/7XT5DuJUxGYBcal1OSN0uu3R/BePxUxihGg5xj50RZGjmva9kLupI4fSfeciJtSysa
bR60LVMkAp7uOBk6msm46lIJzA7htxRifs9lvNIXVf+s+syPSZ5EEz8dr4kuv/rkUVpKYVjzMZJY
qkFrOvdR0JDQhlPZmWBD/n1XSM+Jb5OF0t/0l05Z0p5QTWd/m5TEfSpwCnjnOWrXE7EcnBnY3Gj1
mso1Mp5z2Y2/r92yZbuDjoH+TMqkxgbEohx/Mui3XZ+JUsFSlu6DOLVQWOYK1yC+8G4n9BGF5HhI
4ADBTxJtq62WAeiiOR2FdjnQI5wigfSC8chIUrqG7fyI64ahCcrXbCpLeccfjA5sR5IANGFpbekt
7IsmqSyu96BnehLCtUTKR3PBWwTthoIOxZZLB5qysTzvan/7u8ZZxGFtypTjdYatCdvJNSRqXPpA
Ug5S7V7XxiGHNMox+Tqy/MuGjR4+9Hh+Vph2wLtznS5uOntl0/Ckfc/7xhF651AxEMTjsL2S75Jx
SB6qKw4eOkt6m3IQX3xiEOypzYet/3WW29eY8BWhAw9mUjfrWBVNvJwWYbi7Cnr+3hDnQMuDU15T
fDXGMQKmQKw1xAnt608bvmc5Oh492SVEbqoOHJpQ2upT4wTSIaSjIyoFDjr/WHNYzGCzJOy7aqMs
HdpxQHQ6cFEfTb8txZk3Itwf7bNq8dWYbYt476ZH9iP7cyM6smPO6s42KNRE1QhATULTlGIiihyn
Xq4S3MJHpt4HthP4nWUm20zeTwwoLCVYRKLz77pyOI0TxZwrdnt4MAn5OTP7fTA4yUt2l+uiRvWj
1xe0wVuY6g5cJr7RcGhRFUfhYQxRbNQNTR88rM/WddR863BVJBqOixTWgYHQVtokzVxQYfobwSS4
IawpaWcD9ECHZgP9T+4PTqH6A3qM7c+ghjO8tzXCdrXViSd1lZY2s4WCJhVUZBBP+FIJZu+fMMkF
KNeUXTVLz/yxSmCmu7bkLfm7Ne3AJwZzWoVFvWRzlMfg9vxDiH+bjHoq6MaNbeELryWKU+soXWBK
el6THPCiEj5fUmUh/uwSzawxCkxDg0zE9LRZZ3Fri/TtD2TzlkshRLhRQ1NI+p66x7LFTWogDgUZ
Ca0gpTuDH/hWuQR2c0TzSGk+nLpRl9c/1Pk0Y9/GDMlkoQQ5SAkHlLEkrnbPLHoqkmeOjnPcyrL+
aYIBk7+5QfLRuASmkCRV4eDYGqQse6lnmAaDZwBLAmIQ0M/6PmajFgn9A/hLMOp3EyBVwWRjPE+n
FCPHz7sKMUL8uTW7/hCx3Y9g1TTZtMQ1S5ypY+XKTOoMbmMa/Yrlh+jf3v2/0Mt9DyS4JfBgYW5G
jQ3EA4/kprTh9cGjpD4rIYEjrR5wvnFcXBjUSon8fcqL9Ap82ozCbriaTriBALNevbYavaTlrRlw
gd3mTlHjcMe6Xnv5Y3ct/uOi/jVuOFYCkq5pUeWSWt+5L6/KgCI9GgGZKjj5v7SrLdf25Fp/B4hT
1fI8wDfb3Ly0fQ+EUth5Gfc4Q6+ddFsg4aJUxuz30tS4S9tVt+TVQPCkNRT8SRaGCtzdWzr5s44g
fYydCvgwF6sE2tFAv6AYLHnSa7f1AevGfRWutOD4+wgc4PSR5xfkm5+S6FS4OpxUhA/3kB0TQbAc
okr2c0gK5xAZ2IR4tXF+FY4jBYR4RRrOe/tQ1gC0jAg4LUdvwmNx4bFSn/4RURkwXQ74u/k0zEGG
PaDDFZzSZcq0kc1FFj8UC0rZaKlNY/Lpr87kFWDVogKFPBBn1pY66eOUqPiuhhDy9PBgVkoinNM7
qXbh5Ms5PsBc0/toBw+gFzKyMNkTePsfQ6XivUOCZEcDsQo/gk02rirEXe2ggf3n/IXi2Um2wz0b
np3ey9/fFukNXXLmJ7UuAdj1OPgwdPTCjMdwi6dkoxbV+zNVvminJEKfs8c4uPDH4AL0v3Xzg6W8
aEjGxdAnmvO0JDjeFHyIXvK1VAABIoiJvfeHoxsmzT+wNlKw0Tnb3F6O5LPequ9p/Y4fRGAWBwjm
KIcPsc3bSb8wswZUT2XWnTUG+4wsTFDqpDt+TsReylZy19CKXxDafdB1WCYglTFaj4tnLkQOEOp9
22hkqf2bhNBZDNptJnrOdKy5ixY3yYyjV3PUty6Rfo5bQMOFPhtBh3YcGE+78fbA4LMPXHHXzrBP
HsZv/46qvJYdZrKPgGp6YhlmWdGmo1n3JOFj6ZDZBgdo0sGYKKp5QEHkhTWM9S88vRvLO4lEE84o
ayZKZeHFD43oqiXRJIZI/b+KJySwJ4WCoJruYAtwJelr20xFVEw8FD+4C4UXB7eY4mwzfuu1DJkN
nP7ByulOiPxHyHjPrAe8GGNK3kCapEUJVyJXxVvUf5voWxkinyn8pZM+o8H7FWRRm8+Lp53Sth/b
HHSvSBTIFwnlIY2KxHNyds80qtP8KekhZy3NcnBZZsHoeMrB0c75i6OnzJEmjU0DB93KP5mFCb+O
gHFJt/wz66P1+pqVqI1WkMsgqCjRbNUJIVKKXwqqPAKsu+HFpjVvv8pED0EZPV6Qfy0EQ3txwf8s
zDtIdYANlkdK4xrF8UlO54ioY+zsI2/hJjIPWn7rD3gU6p1S09SBrwp+2akI8jSWm7k4vLROFuEs
o3/gW00LJoRNmaNiSCXW9RY0u7HIdClWgu3Y6ajK2eyALuYzbg+Os0zkU6us6bAE4b9Ux1x60rsR
FIUr6U2I9wGHuavy/ktRYIPBVZP2bYw3QmS84irRSjHTnysyaGpuu7Es1SXq/joa6Lyj0/lPHHud
E8ZCOMPL0y48j7aXO35CEiIwQl5MSbsS7apcbilqAXxkiGdlw79yZpIubNFtQC6jQozDsU1V5usH
alm47F7DrjMqLEcuVV9HG3JbiXoRA7MDWtMKkxGzjmetZ1AeJKSTPFBwxfY3Me/qzH/L07AiEg4a
AkqEAuYKCZWQxlv8fKLHsAaA3MuTbgkGAO/+VQ6LklNYD3zE5hY4+x4bLaOgam5JPhPC8A6Q5Pll
eG1mcT6Q5+XCS59TSFetymJnc2PAoMdEwS3P3bS+EeAInoXvnRLcFy83CgqoBqPljK4ONhXFv/mu
ag8TtDNYr69eWlKVs1w4QfJUpPgZP9Ppbors+DD0y/8wKeYAu+Xy9uUvEWFEtzUlL0KYgBflyrFO
ztmOFnL2NkL03g0nxPCcA5pc1t3a6meFARs6B7nbnbnAYDy2L6y2zWAQ2jmQo7ZQ4dGitveXvrkV
nO1bg6zlBxPAdTmR99/Q/hHg2T16UMSgJpYzBEKOIWap9600obiJa+cx8DvxI3bkPCKxpTZudwAi
kQ8Ou16QT+2Bopdd1sX5EHpl09eVK1EyoCi+9FtuOTX/582e0PaicJAZILNajluXJDrrdKNsku40
8OE5j2skXYlodWiSmLKcPhrUrR6WuhFpbipWRggy3Q7xRKK7/YBMMZKsPdbBNVBFc2ZBtHC5zB/H
4/sgXuFUybwJIcRZmLAhSvmQsBGXCOpYJsm6tMjqENJlsLF1D5dkGMJ2ojlR+qRAqMJkpQ4166hY
IpWYeeKvDqIyqZ4/VxLYmoAVueOOhVgak6OZn4tgVBTmcIlHpv7IOuLiblZ4oY1Gu5Mfp4OPyNlM
kCxcBrdlHJqfvYLYWIQXaoTltltFW00ZT+htJSEa5sGJvRz3ebL/ee7ZHqkyvp7JIqxz/1G9KwDv
+YxQI5TpUZ/ZXds/W6Uqs02BBTZ4QOWtOaVEfw4WOX7oXH5IqzPkRYiUqzJs4swisXtRmxmwKiEy
dof5PmQ9QRgjvOInxyMj15rrpXkQqV85vzI5r1lUmtb+v2mkJT51GX2bEiaQ8SysuLJhlhDGbP3S
DPvqtAeREo+SozAxZFL7/x2+isU6A41zgUpu0SdUlKsU9Y0S507WbHJ72WHxTy9twmu8zSQbfLsT
Ym1ttgqBRyYpGiJO5pAxCrOhq51iCDpyB9qGKQge4E+40K+xfDHxA0WHXEortQmFvmjze1w51BGH
8EiW40Z1i2YgQlFRy7zPXUbe1G/R4TyhnmAY0Yjrha+zgoAFeDoJM8OyIIlmjo0SW5wqUNhCOjrb
msR3mq7l1pWStAwgGjSQTZtiEFQemmPlvMXv144jtFm9Lz4gMWP3GMmwDd2fofZlw55AjBOkqGcG
r1aH63qSiWFbsk/G2D4s9qpnI4Tlx6hIx0SwTyr+9A2IMOTY/FAO7NFgrgih6XucAW9e4OY3uU38
SxD5eYDre5M3H4ffxGTN4sUdZVZcISYJrrz42sJ8kwdyv7gRF2o9Us/EcLLm7c+map9D4/Fgs07V
IMtAns7v3KgLEWdyU3HvhTMyspfSt/3iU8+51nWwy2N7VRW34d3d7foD30U+et02DMRt8uDrEvs9
m1Tr8kLQaYZfUHDfrLgVG2oX3iu6R3kkjemfYXngDSudsiI1fMEnoHXb8buVxQ502grLBsM4AJ3I
IrXNaznQIMCuUj8MkToQMSX7Db9Eebtn+ouRRex12q8Ke3oXORqkqAsoOHlkqN9Olg6rVM2nFEg6
jBtn9dSmGsMpq/TO/sZs2DWIbTDztsYWbkWcgJyydOF1z1zhDF/hYyK5VcapWMU0twrd+Cvnthnn
6p43z83Hui+cRLAv9RdU+T8Sl6XcNCy8CnPrIiDOS7bT+/M/kTtFq6W7ZNjl0LAEz0mAEgqT/8N+
L6pwrGSNmxDohASg4o3o4SEskm9ebZ4T0m0gaUkmvn8AMwDhFa4FbxhuQwg0th9jha9b/Vl1Pd57
iJRPRwd/ojH8ysSsHb9YLUkoOc6TKd3g0HEgtWrsAILadcHfR9PjLX/eNyHjwoNjPWy21cS8e9in
RLBl2/cicokNLLBZKAx4MGYeTfvjrbYXSXBYAmOINxJrJ7af69gjydqGU7Gln+0QR8CN+gz56gOo
pvqV31beHPlmRq1hU1zN1Il7PGMqm9tTqEnEZIPR+eK6hXpsGpO/5J1KQnAvZzMV/fdz0gpAmb8O
QTy/8M6vXIbg8+wA66ThDbX4rx+aGxYeC9zxqtu4BcdrTlPJ/qisawHrRYudH+4R231lNakwmjWY
hyyi/QegjA+Qj2yvsPaGoF0e6cHPM3AkYRw7p9vu0YF3GE0qcL7V3n+u92oJ1bEIZ8TKMfPcLIEH
1M21kdpMFngcC08KSvmb4ooFktiOR+7jhcbM45rCrwYSG/0TXp38rUZ6o1wGKyUEzYLmZNZf5Gxf
7HDbcJ5X9gx6navCWCcjgth0HCtdfUyWFdt/E6lYujx96W9F4r7p/yRcWZH70RWJSRvEboJiFQtS
9CQPChixbNbbJ/+i+8p+rIptBmYghAliQCqtQabbXoSRcn2kNkUJkwlGBIIuTUq4x47Pgnpx7UA7
l1ZTECC1Wa+tEg1r9mAPDJE5aak3TFXWvbzQ7HdzL+hu4yGYQKJs+h1sVDz5bXDswhVC47YgZUla
bzsyIWP001vVq7F7AbbjWwsHMFYanhjo+zTWMFBi5LSNvHqdb2RacP8MU5EbDC5d7MR9SXtY0n4y
z8Ee9uiHpHZPS2dVywshZPaXQZWQaTbHELuNZ2Gq7uZ6sGKFhY9akAIDtLryM6MAiiARfsakiC5u
Y5x/qNFkrWUgDAPAw7qYPkfHuQiZaRl2xTuZhBetrjLLwU5dJPszh3dt26up0y8kv9XuUw9juKdO
iZaWuCfUJQGQckSt6PvOjkFJtFQrFCCINXJykjHsN5o1TjxUKFNSZYrqbL4x1/D4f+MPlStHXkIb
jiA90cYBtdNoMblsLveqvw2i5r+WUJPY8gP0fQQLo8o0oF+IFU7JbQGO/VgTVwxoJgjf4VUD8sbV
p+SbW1bnF4bKWgmZINUtp8TE1RXlaH8P0FI+1keSoiyuFc/3M4iUaJ9EaZBm7zKIeGdU90inlJEQ
hjVn7WlVbTP7KI2NFV7woDAnXM6L9z10AV7OAbbNtJdqRR+Qs+pXsLf01YG/IqBJqx/muOw9tyan
POiu9ehwlIIvHTjE0jjCoFpOTw7NzssL9i1zIjRRJDRGnLfyq2WSJ34EXyPCjbrGKjtooJBGcpqy
we7xmOQySFVuCaEqX9pB5ep7nx1kNqNUwcEljV2WF0qG92BjguLWyBSKnH4s7GrGudn3RyJYIh8O
oyI+IO5gc232H8GC0/rM1BzOkhE7H0W1k9ui3VLJPg7W301Z5PwoNEvYV6tqA5QZcL0rt/apiIeV
FDi6bjeKE2cYtKCA/Fi8QUj1qFLWk8MiXW7y6cWSrniCUJsJ5Orjdud1YI/xXFynQnvHDtQdVcC/
tQe+4B56OHUrQyQUUjVC1w7TVsLNBdz6/wPdSBTtgk8zuLNQwQmiE02XgZyMRSLRzJQ7JSClKs3T
b9YVq9O5tmiSiMIQmCwwKUmg/0ZBNl+B13LFlq5uSd76BkLTLBfFxWBkxWs+1JXoAkbXNErcLfmg
jIzrtHRMsbhlXyadidUo8B3GzFqNf9UlLQ25c5fAcNxScYWk3LyE5pWvKYKAZ94AbzTn/EkwEvCr
IBNIldlqJOORTytq0j5Cf1hM4kRlEMo/pL5L0bbHocO79cK7JjbduqkZIda38tI4h0dl98r43Ke8
yT1Myfgl47g5kPpPvKQECyKuXeYi6zvz+7rMUgArrZkoapZ2S3H7W49KcYtLO2Sw49kVnQcCA82b
sLDgJYpA2t+JjADD1s8TXRBqUhEzSXTQE4S4R0cvhkVYhJhnlyh0hUexfSw7/5wIcg1teOguB6dj
TZzuZM+YNbAsgMZ/l9SQexeWEEIdQ6nTu5QgVI+ACQAJJeBblen5he4KNcIxKDP9INJVItKKhbOF
xoICsuCDJoGubWNJLTptVFrVPh9qguPA0eUatja1hadscpvCdhzJi3vY5erdKj/X8sqVQtkitEeP
gB6q7OHVBQ9mCc4BdqPZNCgP9uH4mda49ubgxGLMocDd3gS7F72RwqR9CUN0W+2GSbNrrnMFYihY
XUkNVNqBNQECp6OMpN/t9CgijoXl9NhuJywQtDG7Sfw83Ktb0fQ4knf0M3w1iBdalRSS+hb1Kf5A
Yt3sv1WFGNl35461cIO6fVAnd2heJEAMPUovmThTmuE4mZcjjqL0zITyHtddlm6XgxSwvbZpW2eK
k1vFLAMNSdxceV9XxsgHTf7htT8dh37Wq0hGRwJd0LVf/CK2awyZ2cDYXZNGEAR3FVH2vwYB4kDB
wQKB5ASKoy4lInazHAN9aZ3jcwBq+GKaY3GrvLgYz8h6PaPEb4blIXCbGtNl1KZn6xM8VsWsfrcd
eNa74FFFyiaw22DZZHFGvazQernyWsy1okssDXT6xoqWM4r+i9q+gnQk2DSOZJ+NMilmDepErKkG
mjJBCwhJWhRLDDuToWzcpL1PKDgkJpwSJiA+wP+0riMps3p+o3VgppDN+ZIRNEGM4SCs7ng51Jdw
OyId6aU4FJHnGbAbohRqmeYMgRnktOB+fLNlVVrujDQmZ89lmrtqfDZ2d4BpdvZfAwXk6R+kXHep
Z3g8Hs5jmHLTuMjdRZsiTF6wkAiqgPn7Vqyk0OZWXUWUJy4vcCFiiiyiwieyBkR+aXyI0sXT2wis
5dHsiixlnknMQc2hyDA3yThcPZ98z+ms+yQ1nduvqwgGW8sM8GsaatbwB1ZlTp0eUXkG7PImqF8+
tn9KsQc7as9CRiOdo+scUh8TOGbibgA6ah9i/5S5+lhNmz6C6UJ11T8YmTo6s3V5AV1HxvMDHWRJ
2Mluqr0xpan2OmE3IIGiPhfBaoUkiKYBxNCXU8tMqdWvKsUW7NubBxqp8AyUMCJ2tEr6HMvOdPg0
Cc30Q9K1WKLtC/H+E23Q2V1+OK85D9QZ9kubKQAS5IufcjQtHgJKcgAAhB2c0vFBeiysfzMfTgtF
TleXEPshji1WlId9p4KrKXsAzs2Nk2dxoxHMLQLauhGXAGggRAJClJYLpWRan9nu4yWPlBqptTcU
yv9Zie0v4XqjVMaQL7LWnFJSwamboJCrUz5zs6nSAgMT5do7HV39jc8I/778E0I+m06rSGDYBqty
ajwKc9atKWymmwYCs0/oHiUmmRCQHrPDQYQaxNde7nmB8X9fmbLMK86uBKBDOS9Wfil6/ua8GVcc
WsaVBsbUjU/wJ/HiJ/oNqnKDAC1oaIUkveuaR34C5+JyEOWoqfmveiwvDpGzyn3gjJIqmAB1vf0A
A//JbiYAQyXocRib83duHjqMm/suQ+P18WUvlks+LQUWQdFhWCu5S3nvhaz6x7i4G0y7Eqautn/A
/7YVR7lnygIhTpXuYCvrIADqYVdRCLmThjCldJy2G5zcPkGwKGuIQ1IzxgxReqI4LGgcJNxv7Fh+
CP+ODLpBOfdU7JskVod8tyb1lfA/yyy6e11FZxaMq/XHEmVP4eDwxxrI0VMmcedlw6LBZ8gBhsbx
C/IoJeDwqL1yRWaTxVNUgqWhQdcBMSOIF/zi9rIYWvxSXom6KRRv7FK1ldCNq+jcDAXgjsMX5tV+
gXoZszgGQcIhtBQrWICXAUUe4AV3WbJmOWMxBrtdLc/rezeD7qQrctNg5Kt8X9VH43P9U/e9fIvE
DdejUDD1QGw8R0icZv/nLZB4v50j5c0GwwdONssr/YqFXQW/3XQPY9uxFzY5GM1SOvdF3AVOZhoZ
zdPIFlHWLb1HQ+5P1evlnWgYipF4ErEQ8zabngxiwmkkNNrPQ/8WfhGYUB8KYXc+aSQrKXOmeGOS
WmjH+CYyZOhC7+Y1V3sRphrTniRsN9BsjTG/yMr5idaGovkZSXxQ/8sihuZ1F83ebF3Ds8A8vLyQ
g4mZ7fUvEmFbs1fjKT9fOAF6OmVTy9DBPkow7ebzI42nM0SoCk5YpkIWXWk04r6pPHonPAtyDY65
hc3kVh2mNAd9DfsW7SdjZHQha3xwBFsBaW3udd9/E7A+QcKxGy/MZn9hbLSBCwdaThxxojFE2phG
oX8LJ6ZqDEGcjbQXsz7V4gmCDeR3wXVHQsdGHdIVtSnzQ8ngFsJFGuYCFrgUJOKo4/KkMnwmA+Re
dsNq3NlJJewi5/mw7EWvrb7SeRaSm4PervLb/M1Ixf6+FSuvmMGlecT2IgnPkU1CrJZ4MYwBsbAi
vlTXsjrcj0TTIErcvQP5G9wU05SZw6kohDjcVqmWkLmoMVOMwNXN2ySyLavgukjRwDbufyA+m0Fq
DYzPxDt95uv9xZ8fed4bQPxPBfLom5XXIquxzk8kZpcnxwEb4gzY62ufKcMHAsFt0vKyw4u39PSS
ZXWxJbQU+2KPkfunaVFGQyG6wxcTOyHCFpDkBv1zxTW76TSv6q2DTKWGOha4BMUeQ6e/5BLOy/S+
teQNU+4Ar2GEl7gpbU6yYfpeLh/bLHO47er9DMkNsGGAKOsMmjAQYpuxZkgvpL5Iq3BUN/OrukjX
p1tMzHybexg4zaFyOg7jTjGVT3c6kEmh8smWT5Z/Z6Oml7I6f47sxvn6iDuAGY/hh9zYDicDU8A0
MTyDX3IAojtwh+qiPP5wO6Wbd5B3IEgJD9pZznsvT6GdwY8bxXu6HBXs9u2h3x5GOxlfVfJGXkQK
w7UiLcANDyagfvkPGSp2hm5D+wIvlM+3oa3ZIPFmteb6Q1Rx7IPGHNypIDb0VdS5sWAZfp4+xZFd
Pki/XDNzS1lvQY8JTR5irQK8mEYZG7M1rq4JeCxE2/V9RBKGOAfV+i1Is45dD/Br7K3JEtAnhU3g
kvaVi+okt7kBLZ++CenLy4/wWtJwffc+FiOjq6xV863ItegRYn0L/zgXlgaCHSiTDFPCuxphZqQ7
SBUYt76FD6bTCZaQYUjVHVkekNZ9+PTWdiodz4uYs4NEAIyDXB6phMhSubRXEfHzmul65PGTpeD5
tO4lIuER18URgPTJ+PkkuDInsGnCDf82XC7GuBUvLM78vFpt8sgTxctAKpXktHVMFJ3bJpAs9E1k
muQJeu7DFMtBZLaHcXDanwOsPEnopI5a1PgC1TuX2l0vUotU2efYxZqk/DFP0dO5nhzOdOv5hZEm
owJpIynqGSCRgUugm0fpLVkmBTY1cNvKhuJVwy/m8NXft8fm43igEAjd5e2j9jVT+NHxlTASbR+z
A5oTtnd4b4aoC1dYADVZuWtlJLryrvmm8FCda4E55Z/h6KLyQLy1clKTjm0C3DI5ES4DZ9YbsW9d
PC4ZDH2j1TX5LuV/RiuS0BGD5k5cGBT7Ob876f850J4NGRRMwgorgvya8DHdr3Cg/ZCPq1j5aK8o
oqThLBmsjt09e2b9aIpf/AIir+qSepkb/T16fFDiM9Cgh4OndcAlI2erj+AUnirgVBskNCgVE/fX
KT9kMZ4ZZBES/c020/+xU4KMpShiz1dP2fPFKZ2g8K2kWr+P2zzhb4tQBy+o1pzuuVz7ycU5/vnt
+nmzIPZzECi4imITjhmlM3V8d8eMtqnHeaafgh83ZUKYKT9x4NS+vH0D9P/KjbsB0wLRxoTgVlGr
YBGriAsbi0AzA+u77wfbfZrQBn2uRWIi4NiNYnlOmo6DxbQ7vbVP1Y6i+JXuAKGsAMr7M5dd36r8
yTQbQCfuK4caR954FOjZvwgUGZvWuQUlFGiDIQuTZ143LgpIV1nH4cej8ridp50/EZaLbrJKFihp
cYoaQcfoFuyJcR16OkvLzIsOtwJ36TiA33lVskKXV+PGk61vsuSMf70g5cu0m2w+mSjuKiCbgxxG
OxSmaZGUA4Ys5f5eIioDh73DPhH2gdVqNjPcxluCua7jO7UcAzmedRrZNEtl1SwJLhFOS+x139nx
6gSx3+m9FEfaoy5gjfZLyCvneB6FI8WqPXZJIFdORBn1oqFNDajau83qm+dvXbwZ0fRLtFNghPJo
9+e3MYdlO2ktHnjiTMNnKRulVkTh6Am1oUeEiBnW05U2s+SdR5GfB4RuGrv7B6rB05i6T/+hl54N
O4KOaZ1v5rMw8kOuL8twV0Yb5+PUvCJglCBOFQ1dWmpFAQlwqkMOHnFezDKbgDyYmGoNDUgTp/9B
OgSJzlrLujS/xT9RYcSvS22gbQr4JwfHshNwgH7O9ON502jods7Kw31NFvxR3Q6fatL9vGsth1l/
XO36oigm3SurGcU6PON887CFgt6eqqC8Y/MUlI2JtLENbaOZDKX/91i/fKy0l4ekje+5c5Ib3aLK
DgSW0RgmJMxRPsxnnfr39DS+doHRCfdpPKoVvOkEMarWnpg3F7pZ5r5zhejajMX491g7SD1Xnjy7
syPSc/z3iz9eFEJqrvzKMO6nJRMGs4pjW07aP0ZRMu8uZ7yCC9hIGfTl52DDZEt9Gc5y97SORBBc
DJHvC//fazPur+I+NaTE5Qlb8RZvAKxsbx83zHD9fk4/due2dUYX3lOXeKGyFoog+hGkfAaGrDUz
T6dMXTslQpk+cpaOAqgUNiq6gEn0KoOYoN1i105qpsMqJPKRmX8RaUoht7j9MQ6wxTSuX1NsXqUh
BxYmMah3mUP4wRCzELGj2XuqK+di8djeyZjYgb/FOCfQjarA9ezNS8MZS7guPyZOE2dSEzGXKzjU
Xp/2mAEJdBnbkn7chD98zS8PWREZto/qXJRSrnV3MBlAFDtUyCyuiRjafGknB1sH/R8PGBtfO0fW
fImxi4ELQKSLIdPRbsIHrlI0M3z1sWaMhTdJxOEPYspVBH3Hw9hR059YrVBkr42Li6kEZHZ9bRSj
wLNKSWL6CWRxDBxPlLZWm3g0XTFfgLOqRZxwt+WvFd80+TsQ9JIEYpUsW3LHYW7261xPTheMw+IM
3voazgzyqX4ANClMz+ZF68JOilGRehYWsEBU0iemrd8fcaLPTf3gnNSJwuwOACcc5Mc8I1qYh71s
41KkLrs72I2/avEcyPbRU8uGuXLMsgCB+r9/ZYwNDpT05xMQFKeQx/EMIoL7cPLgWPZZ4LQpdDyQ
n11BUpJDUpH7gTPjXqUb8axutMGNAa9D/7v0YSrNGTDd1DaYD2s4Qm6HH3Y+cAk8Pb3tHKsAB/U4
zkO0Ya1yOQj1aVi49nQ5Qi3Y5NtJswPtcRCWGg5v4f8oRNfNDLBGjJUVrQ63R/tJpJzwDcV9YRy2
qv/dqhnoZLXRKiAcPSnvSdodEqnx0m+uZB6j/GcoTQwfY6SwB0ej4JyqgRD6lw2HLwDWn+LRiTF4
hOxFN/z7TiI/JJrE31jfqOODENg6WB7sGD2ESYOXzo29ntlQARogo3gf1jgu1Mhe3nt3TURDQCp3
csy6Lh9GuvUDH90CST3uG4D1fZ9aygbGlahdy68q8aSOENv7EI6GxZLpkO90CZ9Ueg+Yxtod+NXY
vqz9umtW1kSVqK7jISUx73kBuuF61Bo81ZUJK3d1n+hJIz/uSdLPe0z6ka9/jQuHWsFSPh3o6C3l
z1geLc8xlHoz7zQ1/Gf0SwG/NDKkd9DJi6VGUkFtVenJPeu/vuM60+tJDu7lQNder19wZA0ZQvbS
DBV4OL9Bzc5UKu5zhZBEbX2JQhr6SVso1LxwdXXBD4DhTkStsSaypC7Z4EfEIzLKaHfqmq6SVUb/
J0O57OXleO3m8v6LYPCyKfpovPYuUc33HSv5LgpAH6vx/gTA0UPyCtiQ2GW71IS5CoSLDy9dvYMJ
sqFsjhVbfba6EDaNSG4k9gfdHyZwtUYlVtnMXdBAAkRqdRl1qRF0GjAIDued+vohadBKIib5cNEx
uH7mDVEi16UdWeNP4ULLSwA2npWKSMwIt6NGzbyDFYmbpcQs9tLO3HRtOMwnuROC2UVjdunS7SSC
7GL9r+ngJCaEReqaJ0m6LeF54i7HrON6FqVbQZpp+xM2L5ZG1a0Ty1a95BOxbaTgD4X0N7BadxC0
sjV25oSazBomeAWaaEg054K5ClgDUF9HWDSu+cgB1RPq6kuC5r5NSlcj2CSACwY+1nmqYQm5AxQB
ZS0CaBZyzdeCYa23oQgC3kAwrHBT0R3aCenznLV4N5tBdaQ1XG7BrBtUFfUv1Uw33bvUfKqUf6JN
SFFXdcYTZ+TN5iRYKwkFQ2QIMnuoWm/2UwMLXYQjZrH47hGHp8MQI+z4MjOChAMDU619AvJwtlq6
7x3pP8nZqfDgp5HT5F9FtsYJuDHqZYPbmHb1kUcqCvG5xynBjnuo7wrriRSEYt5euEKHFo43VRxo
A4HWCOIwmkAmsLWdBkJo+UE0XJsvn6WVs5TWzDcms2GCwXUvVr8tHGIEw6fqNXXZjEFlidz2L3vl
FM6p4YFnjjamlRUinZt39uYZA19sAxicg34DVXOKBWNIDD+5n+cGskyRCEg0PD2wy7eBWDMkCzGM
70LWQecv3u3yeEDvD035qOfp7ndbzVG4kRz8YOawHLE9d18JnpudiP6FU7YBBR6+jMmaZfDzwheZ
/ghwty1EAQfqCFH4g9RzcpG8chscloS5e2vIkmEQOCWDnKnFeCxWtmJ7YXw2FuLkUDoG5PcpYwV7
lB5I+Z7LV5izwNOtqanwbOXkV64z4V2/MJdnRMc8gXtYqvpBopXpnCdlSS8CSgTDYpTNkQsYr1Xt
+WXX5kGvoH9eI1QogWrGzo4GecZ8hsQo65cUZaT444UdFjGuJTbn2wZUWl+F8rqLvUO1Ti2TTadp
tcGX63iu96Mp9BUwhHadzzvmbY6eteqYrneHHOTuGpsRVocGP3rpTRaEkyEiQmYAjSByFrM87Df7
/0L5PgwmN1IQ6H2gioiBJSraSaHqX1qiEU7TNhPLGNWFiEsHSQmKb+o/AvyU+d70ESoZ14SpnPBH
c2TV12h03HeGphfwWRL2JyWJ/BwG0oFOgkLp20iJN4RYQDEs9T+te3cg+bD/sZ2wiLvEweMp4M7b
qigH2BXeroTr2ujzsMhq2Bo3pu1JzMvzYnaRgrlengiRNFOCwSu22Pf6H7AJf+gQ9gFmFcFyr5Xa
XP4x0cgpdNxzaF/6b+Y7WFEoOBn6l/dUhFyRXtpNpq4vLlcsODwEhECjDWt5mdG0GlFpqc0zGdNe
ASdbvXNbdkQlPasgrZ91vCx3xeOqokgNtAY+b/6KkfsODgckO0pTvCuCooFaOCUahloW7lNGIjYf
ZPNRqd8x3k8onrjVdxZ27m2gmJZ3eatAbaYTsrxNxcuYslhlaUHIJ12wEZunQHQnuVwHsy9uG0RZ
EUtYOhRwIB4Hbm8DD2i9xjXmYneR94SsA37babnovw3u3zIDBHmhkRb2TFY0cFRFdSgAFbdmMKBJ
urP/zJAxEsq17wnXA97YIKueS30R1gVSwJs1XEbcKUju75B1u+/vt/K0jYSSBoYPCxy61Vx2Atnp
eJw73KfJ5RIecySfdcY/cUyUWBnQaxJLlfSIko2MTL+Mf93Br/EzSRgyb42r2GKPB/z/A77HQyMb
MB74kWIeDqtGQoeZXqpoJLNsqeDlthsU29UXOnZpiOiVwXVMXC9F9W87KKvPXz5WPikoKcySdGOb
1FA/blYaisV2NSr27aPhefhCJHIjDOCE6qxKCjXxd4wRPzqwe60KwsgIzFu6qB08DFDtdEWs/jb8
/w5it5DBHpIUBrC9rgvGwpPg693ESzqP3I+oS0meaAk9DZv0amPFACGnGftJSMBuieXCPM+UVW5c
m1IBmDN8XY8OyfHIxVGHtsQAve8olIv538rhWZzuporB5xsTze+3Hjpb02muMbsQbdJA6+yv/QjK
P8sIpH9lMPX8gtcg2gN1v3wXpEHDc3KcRVDgj12t4BndrNRvZ/v7FZP6/plC7ufMfJAz2LdBGV3h
Iemk2Ztb6yEWIAfNGh31ejrdA6ggnzkQumbc234uVIuUbarDUQnLCSCT8ursqs6tWOBS7X4ePpM1
6Ua/R3VvDlpFc1QDSRiNL9KIRjCzaupsrNJ3Wwuk7zDcHwm9GR+J9AtGuqAzxaUj0yQRr3/Twz0n
fVoGpKrBS2slfElVQFLP3saPwsLGYE67YGWZo7nUU2g9eVi+MIRAFu3Pz3SWam/P9isXwqKPTY4t
q6sCCHYkLZftb9XXP2lD1Ahnb5rfFLpCtgTFGrtVGOyuBYBrPSZKglQ36HM1JGuG/yND5uxLqDiw
XozT/eXT6UviIcn/vgMzse4Z5N8lA1NrXk++iR8IK6KFeYdNMYNsx72CUDnVEEqk746wBbrl54Q+
DTnL1EXdr636L/1JjE3xqJaxovQRt05hOqXQqUx2NDbuQGbjYkiFCEVFLV2AxAoBPpxLz+vhMU09
mUIuojGHi1vv09qb5zLnD9TZhuK1qBy7ZmSVYDqdj50XEvC3ftz9spq2JILB56Lt5/9WuAukH0dg
pLeVhjtw2+arlfpBlqPhYoN8JX7YekoC/iKwkrxP08cONIhkPFkF0RjALl7wVBDkv9+er8xMw/WE
Bky2fhXytjyllPUH9estq/sFX1W3C7/QTRqXod2IiCW14r0Fe31aJ5gIqERqj3YufRHXzzEizjqt
g7nOYybOWF3Y1x5zQxM0jbDLcbNZVkiOWsTw2jg4OQDRviVtbvi6B/xmVAuLW5tMWJ3JV8K9WKpx
A/Hi46qTisPEZHhZhPe8PEpmUKiIP1D54NUMpTcXlJK8ZXJZyuWxVd06ZqMeBE2hUha1Q4K6yomX
TbPvA7yhassZEpdt5Y1p9KsXw7v3od4orlh1EDJtsGAYlc2cLx2bxocDDEgLla1DdDhxU1VIQZ4R
7EK92J22JzNnRvs9ly1ju/GpSRo8cDWVAfDhKKQdJ4bhIItlY3/JJeXKCsHVQKs2ICO8tYBv8LvG
NPln2RSzatRe8oaneXdWafXg/3U1HXqYAm9tEtKJfbxUrNlnbXr2tupUEm3iQIIOHrMiwxfVrBwy
7HNZSa5gD/2j635XOhlr2t2OikUaQuQUUS68tinO2SSQPW55gLzlrpk/AwKOSE8R6bCQ5BKg5MG2
59CLsTkbTISoiyNI9I8um11hP4qw+tKdD8pw8nxEMY/NRb8iz2uhtLkcnLSaf1oduZIkijjJIQKf
APhi1pBR1gGi5vdhYIsuF40ivIbngWB2I2kmmzvdevTKPGvSeO/ZJll3677q8efg1z7ZD3AjOQOF
hO5cqDWJpYGR9c7ck5RPf6/bhEtmurk5NTppmCtfswnqean7nUI+sqc81Fv5aVj5906w/fBEKAG3
2ztU8uxKqCgshtYfNYGJelhi1UsVtaPyENJmfvWRiDmQtvoWWGqeBO3Tqh/mqtyenNlCFxCV2rKS
8ktGkH7fwURR9R3g3mMfFnR6q6J+m6TmXLCcPnAaVFK59V0BRMkt8vvYZJos43n+83O5TfLKK7gc
VvxnJRxcv8gdFm3c09MEJITJqhBktkeUDwGu9qeBFUQq/2ojTMPmnj8YJPab0B51IWWFUZ3o9PP7
wypvxQNtkfwXTRzoL0sXYTD55iFFeAYcdQrFdOrya4nmaeLQnZ8gnCLjGCq/YR6mqCeJID7mviW3
3NKQmWMOUFWYytFxwecXMqGxu+4x+f2JaWLIdSCV6ltUieWAyqmi8Ln4RmS37LtX0IkD3xPIpVUI
iQLyXOxt/VFCcnO6uAlZ8pz0MnnxCzceZ7BXaeRwwvJwj6cVq7RkGLwlkwiPwUTFPj7mTiuOPjOB
Xdu8zkaVSBekzcmJ3NOzyiR+rIyQzWcJZkfv+aa3T7P3xtfM5G0I8tzZyOkqro2biV5nH9aw9viI
AJ49SweTyF+zJnxW20w7CytGJV8rFInaYlww0Of6O5RgWZgTaAhGVjuAH+cDk7XANjmxuNcutbVs
uVfHnNpbAo4P8aBDtK6jgSv1SL6rfYt6xSGapin0jHt1Ec1rv8d9BGam9AIETYlWr2+S6UsFattA
qF3+9ljw6+Xkczgi1cZVL37i/q5QmALuU2GoNfVZ8gSP7z5RdEELSYH/r/BYR1R7GfDGrbA7TN2b
75BWShbwp4TZstJO6yIN5UyUcPXaqoK/EPf1p0rKfSn5wC5Rtw9lzM9ePAW+6XpZWuv0i0vp8W7Q
khWKDDnUkkySXI5td/aqTSWB30iJ3cHKh0QzeWBPSTYuiZuqXAUT+RA6dLTqvjVneXGgLVKIQO2x
DY2w7k3CeYNpzldzwnJQO6wvaxmfcY0Og2E1EEMYF/HsGEXTFj2TEC6MP6+9Zh2rAdhmxy406USp
ExbKkqFNs0Y+O8O64T4SmSFkC8zFnAOBrBqmbE4qstS5JkzG9xYf4p3JFSiiaCYWrTaWBTec4s7p
evRySiiUmMCxj9pD7GQgR+g/F+UoL/1w/369TDAw9anWs7UyO9EEeDYcyKoBvK42IQIxf1QDDhxK
VJws5h7oiFFq3rK/ESDpTIX560qlukknKoDON/X5ZoP+VbcQnomErVZteEVrszUJs/ZY/Ax9s1yb
6zu6VrZG9XsaPigBy089J6YXmK6LVurYUQ6CHwG/D8BpFdQIkj+9SEevTZK25Y1cqn6177SVKf7o
IZWL7s+lAt172fefVMr4rbztlbM5ubS4f5j9T6T626yXcLlziOFgSDvGvujqBmzkf4gTt1W4/clH
iH6qsrOUDecxEthQJ0NVFAE7wQSXD5ZfxaSM0FdQnvSZLnbkKfLfTAPs4/vYNBMS7JbHhqHgnP4k
HrDevQPinlZb0sKJyoDNEr4VMXLEhnzq2k8O8AmgDNjPKwke29vKg4bvQv9+6Kf6X9bioIgERbtw
xrPhq3q6F7M/pdxyGXFT7tQ9jrEsMmaU50aJjetcVgqYFc6WN0yxvhVpzatD5cKNwk2t4ONcCCyJ
baKPuUJzHsL4+dIYxwGPxtZoXbMrXSQjsRhRYs0vqKPn6BrexbmFslGJrbFMDo8JkaPHAGBr1CNS
yUHPDg62rsIKIwNHUr+oYEv9sDi0HZMomy3tntYlMf5ABqLB7AIcokWgVLclpoZEz1w8RQW/31Kr
Nzk34XsuYBn+b8u4DyvhsHo0cbV8oF88LcrCbMmmV5SLtziVxoKhvT0TjFYib/w63jPs8ja40/SK
KchIbJgCf7x9l9Cq7neSAduhQGiAIaJo3C9leOEq06ZQnU120xag97ytLH+3oW1d89HLceQmWO+o
c6Pc4nn4JSy4UnQYCOv7y9WA63b+zyZd+VQyftKYV12VKka8FLlA9HYPsazdUVU7y1tr5W8P7fhw
TtPoNFA8/CIsEmwsZm1wlp9NgWCPj6xVis8XHkaCuqngXlyxhO0YuwX6XI17uNiAw2lfW0/0EVUG
C3/fHxuEX3lAmPM/hDTF623Z/nmz3s4o1ONdZ8aEPiFFxAQUtFASKoWmQJxcWk/pLXGGhG7gR0Rx
aede25rhiXzN6TSY9kuQIyQVKdC/wF6VcoCYI9LaARF2+rCtvePqDrJXo0lFdGf41YtrRIw8WanR
khRxCYNJ2HRMGo6IvPZv6clHzceKfAVOrAX22uAZCi6JEOqum+4VDDTflea8OksNkZqk4JZwZm9v
qExeCDZkREtM2Jje1Rg+aaACCKWr9CTZtXgErpwG6YTO3wEgLpZD9GlfaFJyCw0hD1N7+hPdl9xd
KbUhs1jLn+8U3TDJfCQTkxckWlk9KF36z+O9fc79KiUwYOpeCG6veFZAGG3kKAwtTaJ9yVLbGtYg
X2S75rcLsaSqLlfTH++pBqcSlc1d7fdV146bRubGTXcoqNB7CqqueMenTzBDAPavBQoFQ/Ks49Pw
LF4Tc3Zl9tRfO/O4oFpeQczHvKIiMDpQBzXcXDdh7yGrG9rJXQZOEeCUxIZG/80VUJ47Q4fjbVMh
7/0XQlS3RCcZxO5WydzwKhuDN7oOlnY75tbdeHvHNz3YmvdTTIiFsTxiymaBavLzKy5Wlb34MjL3
oKD9+EK/vgqDU70yxy0HZu/3kGRpkg4iRSGNM9ksch6dQ/Ly42CdFWmoPkFNYVVjm2Iag7cB8e39
ggpAOqb5xw2gr4JD94FlVaH+KwqQwNC5VRWWtaPnRTOPDprZrGOGRC+KkKipyvxpQoMZawdI2rij
vYGjDfjTsn6cJbV0c+gh17YZ2Lh3j8ToaMwaw5t9BUXGebZuewVs3yUTL0fhmrrkr3m0U8sZ2NuO
2icZEAlMwwDsCSqNtbglbOjO1FgEKnv9PrYM+3Bs5JCajq5LgnoaeicoL5+CK4Oj5QuMOdPftZiB
i1EZlKJJeAlt/dc1wvxrYtx++Ff+uzp9+uMahJLO/38mvp16h9ltHCqALlL84JGdjuXYye0TXZYd
mzLa5hm33Q/vwOJugmqRkCA+JKcid4xL6p75WCwCfgXWMt7kAnHrLhakAqg5LXtB3eW6ojq+1U6U
LnG/hbI3pNeI0CPaDr2Fx1mdSWRrsT+Y+xK0FsoaWSXbSe06MOZV6fT0dCGy9hAh2kbiUBaJ41/9
webR0arTY8a9sAl6oFKm6NkZegGS6nVdC2UMi0s3ObKfbF65opY0qGt1UE9GBXkzmmkTVWCVF4lX
oybeDD12BOw40RXbRJQqr+b8/D985t5nIA6rOzw9SCB7AU/CC7Jplgov8iejAI55UyxqwdxvSi2X
tGv4MChmqWLNZBcPRJOMmUgqibOoiaJTFUDvvqQZjBmgaZJkMn5jTSsjpZd4OGORQ1W2Voro5FFH
sEY1aCOWPvTSQi9V/0S5oepoZLYV5SU87i1b+8DghM7kP4Sl/m+dJxmUO5WybQTk7+aI86M46gsp
UBvl8q1Os5/wVGfU0gvYbQatI0vxc0v5eGAh0Ejq8on0ly6mlER7EiYbq05LRJyh5emts/3amakX
/QyfjBDtfnRC1Wxv1WAZtl3Fjokr+LaZVKt69Mr1E4p6MhjYjbuik5U9P5B2AnrdGsxCgnBiK2ZQ
hfigYvLgKbrdqjO6OlWMpsQEXLMrJaudbBC6djtHiIe317HfoRJiGoFIGWD1IJ1qclhmkImvD+M1
RMicczoA9iqzHSlT2LaAp7CzqGiHFeap6Sehe2WVen0xbY7+qnatdt31NG3hOIeT6+nPqq4SGd+D
hLRM9i48s/iWwWnIJAQIQYEmJ+vKkGoIXoEhCx8dWwpBV6oN/PMNV1C5d8jo7VKXu3M8wtXMEcZ+
G9x3p76LVgjQOvdoAAPPZY9EFU6fRis+MMw9GTqqbuL9q2vfOilRSwmqXtPjnUGp1Pp6qh7t6+hf
yPEE0gu+5Y7ytKGsQqFGD7mwxWfdmcg59cIVXyed/h5wMJVNvFeCECR86QwvKYFgSmxPbf2f1qiG
xcmjz02jKS5mTSd50IkmbarJ6l2qa83P6nc0P6qUX7hfwDeFjNykMKScpLvk2oLqDgDZI8twMLri
/zPVUtwbYu85bvqAeXTACyIMYGtghtYAV30bwG8lAk8/yGBnTet+1dY9I0lazRXEw4fDnxNqHQF/
5v6lp6HYfd80NZt15y/R0R3PS8oHjNwOEhSXhafRZ/biU+Aau1STzTq9ctHGi2iqi2M0GRT7h6RG
K8XIS9pUBoD5qWD9Cbx3ffiepef0unKUfGIYgL6YF/8JT2HBjUSZ+W3WvlG/s09HTd6IEwm0FCt/
HkNPnYx1Izj/9Mmtg5UhlPe2lOFxwVVZBuvRzzkveMyYbvTAAms6+Z9EFhCFxWEjuaz35G//bA/Z
OiIGsXRiSM71Ne3tx8BKvcWGyPPZY6YYIckD+0eMhdkECLPjTLDAY1MnR0/T47EU3MT7MElKDI35
WWwj3HNpANEJIEhnXKvDAh50LL4qKzxeONNJL7977N2JbQduHzAcvf+iqfmeulM8j2H2mn+k+5J/
2Fx37APpXWbhZ2NNYKI8Stc7IJZKAOG9uIHImf+ENvwsYRaC5AcrRH4p9Mqpfd3ZvcKJ3IFZBnRb
wR1BWJ9S91hIklxrU/tsy0Y3y+Xd0gDuSjfq+rymFRgkMZCTK1PUYKAXltkhQt6EZKrOQooxbPWm
S+Ns4TbgBOqqucPH50iLumXbMK6X1nnPm0fF4hWUVzF2NYCycxIXAtYQQflJDhzPkLVhd+5gzVfS
Zu6gAOJ454W63s245tizA6ZPmHK195qf5Y+yWWLGdlLnem3blkajzN3Y1sUEpBRveM3Oxma8rBhh
TkDukMxBlfFromcvI5vLFonbxvDPLVc9nb8cwEzWTutiByfq7ch6tR5OGOJs3QCK6kbECS7V+7ry
iueGVORT2XWVuvwaIv8xEe8gnv5ZB8tFteVefWVd8ZQ9fVxnUKaTxnfDzTOxnZZyM6nA0SLzFuzC
jttNjgad/PFkbPlkCe5lQ5Nde2UmQlzECjuyXQY3yG6ECzpuBbMyZwf0WtkBwifEE+miyiYLZs+m
cZyyXR4csiMkFW0yjm3IeYNYrpCWMe6PpfCtNCr1e7OQ81/a7wA25f9yfdyliIbNEhFsp8iyk3gb
BHCEgVJ3XWJv1Ac23EpoYHwOIf3iGsNnDRuvmIU88izataSaDN2eUp4O6eMObUSDFe8H01tH8OtL
+FlI4AOCHNYiyAUtp+N/kRvPB0ub5P4qxcM8w4Tv1DjRtQmmEWnJiWhR3j/i7hpHIbH6U+2Difg0
yDVSBkku6S26OeMx+xLg76UAvsEl/8hMi2NZnynBcwMD7ZD5sF/2iVQYogBHV432LvlSpkVb0jyf
ezhp3Fv0LE0tbYq7M8XBtooKukkPZ0Z3BnbAPtfvNWdDJmlgCXa3XiW5YbWJlPQA4BPtQ27Hp82J
q2s2XiuMpwOin0kcYRaTLOQzxncPFzIbdPU4M/JTrNbyUyGIhu2DPEKQuQdPnczNBlgARwLgxxW/
C6IrCAcp1DH7pUqLRxqGjNzqkUR4fhpIwOBXsEdpeNiYw4Mpq9etQDgj1lhhwh7Cjx4QRQqqK6Ey
TjGAUr0csk+rffOwCyB42OLJWIckW8Ohmlbf767xFX2uZ2aQjy6+fX2brFT/CIDIYpy1T8JUVglO
fgyRMxUC050WLuRcw3BbweMHx9h4JEzdMj449qrtD+t833hOor4iYMI0ACy/+zViYjkeYDzQPTj6
eyDUv3Mi1SIpsbWG+s5I280n4/N+NS3dbR4jEWTTrGsa0SremmONxM+D6M0YUPyx71GZLpKKGQOt
ZB1FURWgT8NDzdyeisSu6mBMGSlJnIp88Ux6IhziAcDwAyVYCnI00cv+HNQXqLkaIDuCoUIA6hsV
B0N8aEfCH9a+nScf0swIFOo9NitE4V3uX0iYNQ4V9aA1qzBZ9D62/yLBlUL7uInxsNbu+qqvlp5a
fWhEwNPQQ9iD5eg4qNCGYMyw4sU0Z6FEsHcvfXe2nnDbubkejqZacnRPAEGTX8+JwTiqsiQOXeVY
Fj2v9zWlUWit2ghvT32q/7ugcZJWxZ2+N197tjBmM3jcHdh7FKxVQavSyNwYEMFWCMEweKbuBMRb
Fj72Gt90xcOaQ2+9VH6vQg0WhDz+cqhhHZJL4aWwZ2S7smERrlZZjXVzBdeXisf2mEYerZZsCzJr
YCUUfh+r3IFpu1DvzACjpuIqwI/inOE4T0UPn57CoE37QEWtuRM+2sVI2M7uqTi7aWp5gklSSmyJ
XBcxuVSsEks0Ht/pc7imO0u85XShlttYdsCF6uXLQv07jiRSfVfO6+S0Ae96Bl541Zl7ofPRAyXq
FqZA1M0Y4EpAxUFjFUn2lEGZst1yiM/fx2lrKy7kVoG/f1Vs1Ev05hKijwDtfD5NkiQvL+7/QSYH
VenkDiuATuixzme/QYBJ2kodhpGwS2Dd5UA6qztjrlO9ppOAHkTfOjzVsxLtDscwKu95eKGvH8Sr
CRTdYND6YUEKBavPUF690lKWmE+8Qhhz5Pf+r/gZIqoXu+0vMmuEN3oihrH8JM9+yZ0HVqvMjXaa
vvA36Rglrfv2H02GDjSZi3x6bMxWdStcXX30Otpo/9cKYnPlFqvndJShYNUeHFmERsKX7rkJ8TbE
UEDp1S3luFsFyfohNPRZJtczNDcu9FQK2FcKA0tAcypA1F4+q7WCyRjhl6MVrCLNU3/BhkkPFoiH
hRY0uDqR8yhaJvqZklADgvfYgqR9sPOhYVhZt5uTWDfJELmZPPybbihsimss5lyRBko5+hs8C2Y7
+Ls5VbNU96utN3Rnw5pSNnLu5v4FMNdCzCl7FTAo/ZRlcZwRm9JRd1TLMF+KNDXNEgnhALHNrZBv
jYPuphT5gEL7wUEG2QGfqsO4Z9SHCiaeh1V3+vV8+psmxPeGe+euiVK3hOAvhmwwr87GD3s0fpDz
UeoIKdt5fw1OiNOSXR3iEZ3iV4cMThIeAszuugOvL/11MWviAfatKN6ufNm2+n+gXbV4R72jZPCG
itFcig9nIJuZ/X4X77KNK8hDq3mtkJOqOabEstM7lmqKwQtTQusnJhzEQLLG4Ctu52+qGAVe7Kmh
9jgiBV46cKZ1UT2u7z2uYA5CNzy/dD5ScrInKKozmFB6tTSTuAhR/iwOaqpMNUUhBmPF0UCWDwN5
GLIovp4Qs3/6Rl3dVut6C/ZD9yaTDwnMJ/A5NGrCYs+BIs5fdODY99AegFRrqDLfQHBRGJGOC9VT
nwpq1tc6GQTGwLF36hxEA7Kak8TxSAlHkMMj7grtBm/ot2+ZxzvfE/0Eu+a7T4U77U06DyMDXHIL
zDKOd8z7qVq44kXeBWL7FzdyjWmEuQ1hzRUQ/fQIUhzV/9ngqbveDMZe2D2eq6z7yU/313liNFhu
wAk44hIji1k3DupTUJPiNFCf52r/uplTYaO7WV9pXFjynflcoz2ynfgwmadxKszEJS2tU6mAi8s0
M48ArHgXMwuiKVr9HqwEZ9IUGIAXMzss45xsjVKzU4z7jEVqr1HXvt3dRBngo5P7f8Q35JQBtBCR
qAVtr+B4ak0/7MnJESFNUXQAGG4A6G6PhoL15xCgOBDuGr9geydP5MG6nrUDw0Pkj35hmAvGHCq6
ki6ln0/QYmjuechLt4SkySRcVQu4sbMtWfL6C4pGBZMgs8vCEakK1Ah+6GoahOd04Zy690qhHD1W
KWOJdS59mvp6Ty7b2C2RkUulhxUnKLM/N6YhJB+hhM/Gh7vbK99QJEs6udCNDNqry5CuW2lNV77B
A7LBd6ZMGwk8AUML2fKH4b9Jh2pQZyEUTxdtwXbXyORyS8OQHQr3gByLN8Gb3FP/m1duTZZcufQ8
XnAZ1vMrFXzuo7IB0TK68kibGO4x18Ct1BqbAeExfm0dvvk1rFRP+M/4Tti/b/Em6k0chXM/man7
SH9nuzpeRVsE0y0lqJnAiHukqjs64zX8C2K389NRA5kwjhum9evdyGhUVtNap2KguLx/+2VzSmNV
5U3+Y8qLvraUWWcocjG5p17K9B6Fg5qRFRwtBNx9tIm1brO4UlSh5BvLz1GiKnUwTZdIrEXIlEsR
7m/MW3qpoqoMl1AxVh/YzYJqglIDpVNAKX/cMk8m0UptitpR27579LAH+koi6TOvDgsh8A4wVSlC
WDBtRSQNMoZhfynlfNqaYp87dwQBic8pOlLMo6sIKeK5bU0ds09OiGlfTlWQLbxt3aDkDQTeebv8
hZjEuZLym+aly1pClWp9/znelsSSFvVbdRg3OKB3ILP9zTIkAXZaIxpBMUQEZHxaZ6mzITyiVVt/
U7nZYMjse7/lxMwgQGuUoF+EFtH6DjzJLtg4smifPwoTu+o/V6weyUDiG3WvZU1dfK/HFvoDlHrj
N6qF41sUuPXeQ5avw+bsQtJW7doJ+MRDa8fkKFwYzjrABtX4uoTF1LMTFyxWiSScDnocyUK/9i4c
68fXYepwCMj8xZoKN/6iDWo4+eq11t2tlYnwoHyyRUt24ub6zOgyuRuFTdWnOBnOuSItNaLFxf1N
Px4ydrydBu7tXK5J81XmCpa4lbEKIjQikHUH3M24jSBMSD9QYkA4Ro+RR2WffeQfLA775D7L4FUo
uP8TchSjAlH7drfN3jnR4P3YlykgqtCVwIZNrNU4i7xklOQuxRWz4F+10N6uTI/dQM67pozO+vkj
/bcLIiEtAO4ikA3u+wW75bG6cKXogf4MT989wjNJHx8kDmcYfyrE3TIx5QYV0bCL8/rcJA0w9eaP
1Soguv83GzRCv+1R0pXemc81Z+ijblKv8xV0gKZWnN2pSTtmu0xXLY2/+p0sP1Bv9oKKoat7O/wQ
H5mdjR82z6o5YMBeqajmYrkG0yj//XJNiGESI/JRBR7+TufG0czqTuIndCWNnRePA3eumnt6zb4S
hgXBvAOLxgjntmxpLrJe7wiyux9DccE3Sy8KTwDnCowq31Dr2BDWUOIAEiLt5BzvGOMu5n6Q9z6v
iLfm5z2BB9KD9x2fzwgRPmjwqmwfUe8ctJ8kwTJ+vii958Y6oYF17uykW8B3mHlgSCvhynOxMLKs
+Vxt+1t3EenGJ84Vgyu55qAh/u0TLmhjfvf9KqlPS8q7NK9E8VRqrZNrB0+K/a4AC5qsJAM+80vv
bmPzE0JlcPW3dzGcx5FcG6JwLR4JE6zmTrWT9ZuBhZiOgsEqC2BeX5luHuxw0EhsFtHmw1ji2C75
JFdqNVtWzHWRlPJmj/E1dtWmeh2GYMBlMxULOINGXm6X07bYsuK4F2bpJeq2BLi4/M6NuELwaIo9
XKKozhYIPi9IjhVBHqWpZIUZeymXKHXtEKPYkU62uzdCRhwWUyAbqanS1/S6muV08Y03aFQyyMKU
Uaq7QI3jbJPRn1nxhXZul3egEJxiZe0PNDE61JQmDEhEAtuQg4w7o7f+k/f8/3NU11PEJ6iwMtQT
ZUobybMN7jQ4PDqINPcI3Slt7NCGp7jpke8YRnxkC8MzdyZFCWAhMfDhGObXpkl88laIK6Rodyz+
Hzwl7xxPtbrqfDWX4Rq0sz+C5K3e6eAYmjSnxkMjghxJg+68aaUibnkqQJQ0WDdaMrGETCZTATjE
C5dg09139CPIpRgV8jz9KF0rxy/W5vXmt3l1ssGOiwrDPt7XGBKaDyAPkKlpc7GEe0n1yvLWPcnb
GdCAk/zuQbwx6MvnQBtFF/lDmaBMjDhExSjLJ7cRAi64lhuTr9ebRpbPIK+4PENSjTeDLOY0PPFi
3Y22I0unORKSHoK8fmAG+2Jyzz9P7kXIXS+QfsZiKqeVquh0pelpTFTcTvBNKQr58WejvURVNI70
8mUJ5mEHz2OB5vAtYf0z5U8FbVElCpVgJNYpbwdPbKgIWwgmoCDqthdR7GR0pVUH9a9d81zk/I39
v3QSa2GmM8+R+xuJtbpI5RYwbBWOXpXfEBXDmyTmiZnm7Znm8eI7nDmwXknbO6UiKlsoekxP2/4s
7yb7LAbhNBtQl8pNokZEvt8L+LIHKSFZbjCdaZKmYW9KKw9+8Vfxf3YRP/V36AR58hhLmdMSL65p
fGXkHS75g1XAAE17XNR1+r1R8eEukgAWQ2BEWZfJ9IVAVr24Vaw0iwnDbhZbqukV5+oeAVsP7z37
Pi+xDiAoYg1rL+2spGSqTtlXR+NIYFZeLdrQB3wSH4Q7u0Oog0l0XICUHNwP9jLnkz3UF9IQv9J5
N3PrQ/ZYZJuL7wUIzc1Ij2EswvHXGy1l4GQ5KKkmy+7w9wg3Xxr1e+CcpRQQNjh4lrCuA7vobmRw
w4cPaWUzX8l8NcTsrVu5j2dvOTZ6ZcU5hlPiPNKW8BWtFwRj98dlLpxXSJHYNG87q4UotZ5km7mD
xwN2T7a5PxKG/K7abNOOh72pa3+B9XXE2kGAHwhJSZlmQ6tvK09KgJdXvvPIFIGc0XLdolTW2Q9W
KkJQYHBsju31c9/lg+Sp+1ood9I/+gEQuGxiZzB8GhDhzu/bzrsI1xGiG8i1ol1oK9g+lzHPKtkI
8OwvXv+eDKCqvruykkXXiaztyMXzFxUJvuPte4BDs/+PkWOQxYqSWZDobRpH8FYiviREtIwjYk2q
faDUhUjFX3KdzEgVFaBOi6nW8+AWIMtid+0OA428kKAYLX3Dbus3Do4CtdoPEioWu1cvs+pDsAIo
y64z5sLU9LbwB5BWGCHlHgILVRgq2HCAj9XzbqueTD3FE8FT85WDAGhAVEo3f6gnGvkwPPpY8HSS
7Xass5dTAI78wBnrLoCSKWw6Ug8tcbLF7yTE2rDkUWWDJHk3bRyqLjKJEQNhHioGrrUkXbqqp0Ea
jZW6TF3o8aVWUPr1o6a1Dh5E8Zp9bsxctnqpvbaO714HOT0rgX3/6xh6NNkquESRmkL/4pXBgjuk
lkVxZjwF/q1jUjBrVxlobgjEPELjcVSLmmaXlkkxPBnNWkzGM1vZnryujnNpggMn8qAjrkUM1LGC
FuDp1KEmtGBNaRk/IvDaE5VHOqVK86fFZsOTHCSW5kleIfY+mSTHZ81GJGW/RZy+XvUgFalL3PvX
A2NZq4tB/wjU4/4Zo0tKx4K+/TY7+tBt3QQHa70UosaefxfAT5wpaYO/B5RQBqrIVAhHF4tHWVAg
0rgJJ0mZaCiHuA803aZ/SD0lf4naa0/osMvxVni+1iRVXHwddDaeA0ZvjIaOoVvGCgIx9aAK6Tnk
NHtjXJYIYqpRaCihkVRRDOh5R1BicXCoNVggZVzGBq+f8qCZY8iNUuM4N5Q4MS/dEhceacVjurAv
0MJMlSUOEIQVRTXw9WK/xomvkOmu7BbmdkQSqo1LQFuJgNO1Bs4RUVoKtdX0mhURjILQ2AK1JCVS
8jhp2H7n0kJVphg5BLxq4SzfIF4p1JC40QSqwaEJAdztkPpeZxFt4+1xrux3ZRikXpTpuT3jTSX7
o/OEJL0nxfCb5uesG3DWwG3bxGwA69NSxoLjK9esqlCEMHNpn+2XR0OrY4Lrtv6KDsDQmIuJLrpA
g815dYYuh8f+HCkQFTGmu9xm5/kE3MCpqYyk+flzP/y6e4XlWdS4OdgaWyM5HCzpVlzmLqnjbPp2
92PRub7emUhHc4X2f6y88y9q+P2v1sBDMLc5gyOofJwSRp6Gya6V3hHmapiASDwH9mF4aYF9d+wq
k3Ff65GS5D7MxB/TKLetmNr3fXQpNXDwf0xa5TMYawE3nCSiSmgcr5mRyvKx/huTooQN9AW35FwG
25snTlHXysua37yOxQlHukUzNulR1+iMZyh3Sos5CarrppBM9DDXB5Cg67omjLwgj8S31xRkTRXN
vGwkEPbhZm9jZdZGoLfiAtzPTz77KDWq6z/r1KXJnPAxdrlvDabFE7kh0EDq/ePyehz7NHUrRLS3
Uy/TFBxXNBiWw7q6PjMBnMSqrWKG6DTH1tswXOXQU2RvHSy8URv+qkoZ/RMf9fwfjjrJYK16dvI3
J2jpuAS5HdqFMh/qFozEvYta9Y3SJ0CTm6kQcph60hQPSz9yvJLULNeZm3D/76EqWEsa/i/dE0oP
WEOp6hFwG6w333xzzonMu26d8voqEgh6uHmfMtgw/ELDPHPjTsF43EkjxUbd21rLWBu2VIpKc/mx
Im/4Ns4ivFGtuRn+3AJumBd/Jwo+Zvsq4xgr4an1Kol+48w5tfZgIGGz/SgfGcB6SAmhhRoMzs4A
vYm8pXJl1zrgT6os4q7jIG0jbERsszd1k9FQzeIgNwY6yFRPzYKbyquX1+x4ti96z73hQwbRbH4J
VG/YqAXi2Dyv0ebxIx5v9GLIPAcz9181Jm5G8jhdHCFU3MDHXyb4sz72FyQlw4tCCLAWaV0VL1D7
jvVyPSe+b4lu49TSI4zZjzOBZPA3xMNJ3de0S0F4t0YKRmgq7E91sEfKHZ/D4t06/x87Ip8tGPwq
29ehY9DeA83nCaTSpYzhrrJIVVwyCVckkVERo7eoLyUpMqOD4pN1avlMDEhOyNBeb2doBLx8r0CV
ux/+jxDjtwzYq+5MnaNYw7fNX8bRl0htdeCc8EXI44Xg/zH3ppg/WRWBKfot7FmzHRW0xhfWQ1+p
mVeVlVogWIgn3IOFRkxDRU+A5A8LQ2jYPHOyvDJvkLtlB+nBa8Tq74l8BuBS5DXar8iijiFbNKu3
IaToyYgJSPJatZwJdSxCK3Le/EPK4IgxF/xWbzivYHh71BZ6lgkCWKk78latnfFrDJVyzGYUmAjF
YyAV6uaESMgpOzRhUevRJTs/smRgSn1LqEDcoTJmqe9P75Op09oAwB31h6qHFfyeuGu18lm0eJmM
qX6kgRUS5D5HJa3mZ7RkDLx4AvAIR98WvZVtW5kk5yZoUWgvJJZmciZ1AbmbwDvL8g8oxcSBFNGG
/ZYkwJiafShMWDHDqBZhtIht5nJVstdOfBxrcoPeByTHvlQq29WdUpK1cSmwfpFiHX/zqIwNMMoR
qBMm8797oF1wFpPDV3sQXmOCy2idvZ2T02BfVyFre2KAmYvT7lY8aseFkAjRsVFjLhGi9ZeixRJU
1FK33d/WWCAifOEZVHvXbYGyFvdY5a0iD7YjY6hUzaZaOcYfW25cY/cR4zytrTK66dHb9ysUWbrr
1GFoP7pgDzXLt04XB88y79pCg95uaUYhWv8e2/eiWOwT/66zOOQiUgY+MY1Q+MqIuuuuc0qza6Xe
zdOSe4LCrRqEJL4HyN6rmS+IKlLNJ3y11gKERgpSRXbcUfR0RwMDPeWNxRBA3JqpsKat+CtxYapj
4+M3ljRb+kr3Y/otrq2YFdwy/HF9zL1SXs+Gt7LCHkr8oinLzCigyuqmZJ/aWuH1KXSzpvYFvPGM
gV090PJ061dMMZ46J63mwYOXJQ3biBSWOF4/VSTNWxIvplzZQLhhVH54bwerU2gZDJu/2j4pFp3U
3qtZX3qwQLJcIP8VZwfZxgIe17zKVm68LKrhTp1q/mn9hCBCTxpSlXS8k51aaQl3SsauMdbnct38
JMabqyg/q63yWDGrXRpshxnBqqhTp81loaeH0IH4FnOTvsKWwIpyGBOmdDYCgZHh157tYwvN99km
cShq9pMi0oR1jCCEtHoXNZX2SQ42b2kcvzBBSUucPLuoPe42s06mToF73dNaXnSRdMS5WR0toHm1
KH0AiXcJz5n6g1OGsIR+ZG6cwgQA6foYs3feAm218IA0MkqPrpapsyVFYW1TRV50nnAFLnYmkQwW
6xA82u6GOn0/PCQotc7w7k2puYrrkeCxm1E70M0gunUe4seeWYafHFRAG+adX58hTAL4HF2rnndJ
hYBsUcmun0h/BpssxsPFumyA18T/YDm5ZR+e+nLW9KDOfV2FgeSEaFmPf8/PxWwPMLVbR053ECKN
SrQtFCs/UCnXBQpccsOTOwzxC9/uwI2x/w8amLnhQ+K3czeyQSiYCLNujpgivrUF187blMakVKPj
ejG/ryCaupStzxmulPQ35oN2diSZuM6GZnbDtN4QDBhvVyMTveuNiGcbUWJECe7fAn7HLSIQTOMS
B32PcorBpDgOgBGh0kWo/juQMDccDjmCSjfjtKRgmg6Tnod9eezbWDmYmGrvJMMFKsFn5OonYoHI
QuMijL1Hqj6lo8fciML9nFnEZXzlvgtzajPaF6PHMOW/WQcIKwNDdAXIjVnbYrwmgM99v8W2lLMv
pXgotY2z4p6AZQYLReC7s78dvmbUmQJy837+EAHQBMYPOIr0zXG+kmVjruWmmZfql8ezp2TGzgXJ
NXRyC8WOcOuco+Y8bj5zLjOg38YLP0WnqrCpyJw63iseZ29tOZsa+iWLjvLtKnefDcfTajbUvMkZ
JdvJEphYWkHKjWwrUzRhAM+cJZ8b5vt78pgVL1iZCmhH+0j/iPp6YtjmFYpZ6TZMG6xVhgHzUiD+
gF15Vr51greasewz0r62LMDK745EZGqk1a6eSt8KwIT+ObP1TRToneIh4j/RHuGt+LUCI3/F66I0
KLB4lSv2Nu3/vOSNmqh6vwYpUjcCnxhlcjn34kvPW2uK40rRC7X5beqnxH0DoR2OTf36J5QKJ5N7
9BG6dnyfcZIwwSWxWg2QoQ2lUzUyoXfn4G3AVNKpPt3rg9RyFu0nOHCufnKXc6n/jwXZq/Q62CZC
UWJS1d/cf6xyAFChVIkfq4DMmOmAwdtPSTGy/DuB5WiQzFXHwYeNrUPu5WHwFDmw45s1yTW//QUD
51H0Wnx5Bj186ysnaINPxNtnWYqK3bgFdo6FM5sSUjb0q8uafqCMXEaNN0Mt92NOS/LpqYC7/Z77
o2Ay5aGnavtH9YV4QEVXRrNI4Tog5g5b5kez5H+akPFseKpj8sWDfS2T49CGLNoE9H4S1gmkc0S/
btcpm5kARrxUJpV8PFF/i0pP6ZbpQYZH6IHFMDirP7vz3TBR11HiK2XmHOG4Xuix3L5uUg9mSncR
ryH0/TkxobqFAoZGHOENeNsk+XZFkK3jaxt93qJbOkygP7gX6MaBzkqg3OKKWF7P4mSdaIQkvxm4
lqbQFKApq5b7lHZUirqOTBTjyyqTFqnee+rLdef0tEYuAefUG2Az6Mmqk/WuQtceA7M9mVGkpvN4
JzmhyNhXn7Su3znSwy2hY3F/FuVL3eUKsQY7t3Nln6K1X902CLvLkkuT9xlYGE29FcGka/jF7Ej+
7NCafBOl3PmMMNgYijKlg8iJxqETUMNsx0Ygs05N0EGArUJTw7GsMQxfhD53SgLnXW9/P36sH6Gx
AoupkTGkeGSutktmouCTiP0qvvx1bkL8DRaKfdqokitexCi9b5INFiTfgmV37HK86j8DRotfIFH+
wkEh4ahwH5oiw2IF0oyCaI10aHRYnTqxDYsNsQzJhc/KNicetEX1vmy9dwPS9G3qG+swfDTvaiex
bGrrRrbI4kKXpRdcU0RwZ7DW/NVRpyc/9lIcLqUNbo5BOCN2mL66/PQd4uU0U56iOa6nZ0hkymJq
eTvjU26mVrS56dBjQdeosayiNm9BiLZESyC5DR9lrgzYbLQnmKUAX0hp7yGX0GRHcg5S5Zo+tuJV
5tmtnOW0LXCDl7tA9afdz3WJ89jwCsQ1mwcB0tjUjcPC0d1dEvOisMHUKkR3Flzz3/7F+FERGV56
Ph7tVOVql2t65HbaWPpYesmwBIxPPg3weRvWhFu6Q3TPpsHL6MG3w1rhd+kl7CWcYznzxnEEmhbI
EL7RfzxCjbvWP9j5q+0p/MY49VNWpBKyhF9dN1646AvEoNyfpKp2DG6HeApiZpgfccYl3uDEOJHW
LIfNxF9nwXL/ZmMHQuIo1fDiy4jwFvmlpTe9OohtOYuW0IK0Acd4a030WP/tdNInBHNAH/9M7xfZ
nQumminorR3tr37mft/lnYODuZM7u0FmPsbc8u3UNCdc9uolI0arDRiVDh+VJSXmno7q9JFbJiG8
PjqhxE30de4A+vtppUdDUdjbWKZxyholpxM9pknOto1CRVUflua/Z6QbnAESZWoWs59lUjOO1rhl
yPjc+uT0JG44qqU5aILvumPK32p5VdlJJAxh9SkhYyFcYUzoFJNsBUwwAOET1jBD5uA+kV/eGhzr
suJKFZwSsKwjDT9lDyUc4zVCcfPQAxUqaDqDmIuzBPaKlYmjZcwqHN/d+Lwgnoe3iIRpYn0jOA0U
mBXniWcxPwONBbIANlsBdd8jXLLke/almWTSZpETixJUJw7labPNfJh5uTB8j7twW2wEeSuZIz2b
H2Vhf4UwNZTSDi/GxQW7bE/vb52ttrlbcbH22a2pXlETIgTydbymCpt5DjUWGv8GW+jKXJ1rv6yz
/ZCkCDUxZftPgPDfbDCeblpuw5C504aDD9DF0Jt+X6fQn7YLEWX9Hfb/71S32OELdqjdBceXV1at
0yugJSDvU3J4X7SOkDVDu207uo2lDeWZpgFy8dUt6V495lgGp4jB75ndvcrxj02eZNQ0JwhFgiPe
jhLn1cf5x0BA6uf5Ikx96DCLEIGVdTX6UxrG3q3gp+/H12m19IkRCuEt9PKFVB3zzMPG830c3x1i
ORQKN+N8I5Ek60UgG+/1d526ox1FN+/fiMcq04MSw+acPiX0kJ8pi97v0snWLZG8APAWdENnok31
sW84NLMHmHRCjmb4kc4qaU08Vf1naxbxp/H+kdb4aj0406xjPWB/Ymx1gH4M/VfXe/vdtMk5JijT
QgJPknJvfsohmWaIRXxkkusnOvqtQ+B9lP5kO30zWCYQguiWTc9DPK7DZ7KTUgjUB6XxQg7DR/2j
UBdh1ZlzVGFiYooEAybsERAgJ1uzVMTP/iaymoYKHCtScDotYz9t+TgYEZ19zrjzknTRtp1qFQam
bsHyLk5MWIZxu6mZzkAB2lI+xQoXvAasJfZt/QAdHET+2fvGOzH0zKe0ONF9e6yg+P1kB13sOhqe
B27PJhzvQS3UOjTM8Grbue6ukxFDcF70NMyZJ0LrzyXmbl60jmNwIzyIWSjd8ysRDkJjgjTGcung
JC7nH2dtgAQIu9FC6jvH4lAzjTe44+8A39kx7VdE9rQqR7l+cmNdVIeWechMWKNrsB+XOEnL5Ly1
V8mjJ7IE2TgH0nNlD5CGxJ9HH7VcVkC02TmpC/i5/zvKVac8SRO0iWRL9Nfoz5AESF4EpZTRxMRc
PVqsqDyS5sEY5osi04E5+x2ApRQRpO30WE5Bx5Aj6zi5CO6MwMWygii3J4hgr46JaCLzFcO10c6t
Q9rBAOFFmPBWdaor6Xo8sha0pC+KlLAhJMvOLXvoPu99594Q6XwFpZesV7h+pUzdYFEIkORph5/m
HUZ++5XUCAI/ZvzvJ8SuEm6O8TgZkfD1WI81bUtja0xoos1muh10jnVHslxcwn0mM3i+6VfYWpfw
YY/KmHtE31US5BvQy0Y/59j5ZWypbvppFS/MURuC5yTiXD3BCwS/+CaGB5uV3vtZYIozO5ZxNq5I
xP8ep3jf8Cy+SaNWv6MjF4xiBxRPDtTJ5NlX23v29dTHbTdeb+6epwZ8ckI5939+2E1bfmV+f/1A
Un2p1BDOM7GDxQOW7Yt2RdYbfRQ7M+8jGo3sdkbwHOpKtoTvo4Emez0cqmjR/umKSfZzk6PLdJ38
CW8KdiE/uEoU09JhyXTe8digA6QKLy3QQEA3UVRBz5lBZeXjV6o6rIXQxatdKv6xvznPsKtuk0Ak
tmnXVMJpgAneoVM1O+1V2tiwmrPHCgD2ZtwDpYqyOh+7PdVsVb5J+65rKbpX6iW/rKlYlwgHUVZd
sDCsovKF7cefmgjuKdn5V/EXiebXl86NAtfb2YeYAXk3J8SKogNr7/DMxNvFFPCF8kznnBShz5Ws
Ol9hlTlABzTC5YVhuGoHoXTxQ1lFwhTrWnCbGgxu1N3k5FQXvc90mnswdpsUudR7brEOIkO6jSNh
VynapXER0T8VVVxJD9/1r1D/KiAzo0V5VXigjH/LM6yUbpPPd1jkP3K4gMtsN5/RxMmfiKIvjm0p
YxqET4QiDc1da9iFGy8cVNtbrL8Nf0BM5fb2HprROSB0YwJ/rLHg70/hDvIS5LxB47gThbX4tBOG
05J/5SHF0y24Cv/qzUYGrnQ6r9sxk8mweQzc2dz4gfq4bjh+lrSY1nIumCTgJL45XBHwenifgU1t
UQGe4Qkf8GpHLZU4QMRNOLJ6wUWZ3fNEJFwQay6T/65mh7CZzzhYrbFGqTb+hOj9uM/9hR3m46W+
KKLaWeW9gqCKvyL6FyicxnbX6Vl3mbcC8XAp25POoCIFdKHYQ/Sb45hSuJJGMbFcplawwsAhdMqX
9TXMZxcG79b3FN77L341yny5CevYcOy77Lg14XHLXaU2mQUkDLaP7ePmf3WNPaOTU9tKtZzFKLhi
vnH8NyRKjyGDey12A8/g65HCQh9ZlA8OAcpVJ3a5Sdz+o9PROOQwu7VR1jFCZRls024x3dkFaHWT
4y4UxerGrSDAtnktLdYXT7sRwPHNk/94rP5zDihE3GHpcJDxbFayQgvmB+s283cjPZJSP/X0m233
VAnrvMNREL9BSQUlS1ozqSjGudCeYLhwfT02nfmImSlrOQLRC5IxDLpG+Le0zmCfaxV1abitFGEf
+YQ9hNkHBxoENepCK5O5bXQO+Piua2Mevhj3EmRwO2mxUZnpo+2LeifO//fMzuRLuTMyEulWTuwo
i/LhEpEdINpIqZxVy07KIKzl4osZI6cwMAi5AUqNIA2HEdn0rU0KagHk5bVpgOgPm0yQEFZrKu7D
qiM5O9lPl1dAkfdeDFbxsq6eULmJJ3ruIwVVwhH2Qe2M8FR6J5AXzez5BqAOip+nHJkmlooQXeTs
Ru1ctgZTS/6k2zGFgv6rCQ8wGcYB6H40TnhlG5OlhFFmvBW8rirn66mkxyihkx2/oLSZS0UEKGo6
IMJV7dUzz/soTbr0zhp7n1E2pta8hOd5rXtmk8FDRPaVzsV60QEuG7G+U9uzObf5Xj2vqDoZNJbm
tBD7GnVeKNl+GottaZX0NJ8t9sA/eIPJiBMRekmVSpvs4ntLjyrQQurMS8YsCoVJfN/CQrDyymdz
L7lUtwJyFkdS6SeVJcUBbtV4B+Dq8FelJcSKe1a0tohojzgNkgAKWaWeSqhxab6HTga4QpDSMk0c
AOzhJugDAKy++FAPDd1aILnQGc+8e968mhrkDk9Sy+/8RlgTzH+QxAx3PVN0vaAQDSJkzHF/r9xI
jLom5LwbuLaIBSNUw2UKRCUrtSuH1DO3prwQHxJhPIJa0g0yD9WkvbQDDidXD1tClPHMQqeUNBsM
aiQIfAskfgii74sfHy2nYYAE1uh4zinVzge9uJaEEvqeOHlrBwgU3HkS92UN4Rzci+Ak71tjbghi
XiV+owy/Hik+Lsn+42iPvAVO3BaUJYOYelxP3rpdAtiPHISDDFqwjArpz5wSp9mZ/zARVf+Nu3gS
kuY7DKus34sog6HOEojzSVb/K3ekP5GccN6lN8Be/58qQM2vWWzzWX71tYFCn8JgC51r9UhTqTWf
2XrUddcnL1W56OWsa7Yk4DkLN4JNIzhdlFybBoFpaCvrz0yq6GxXj6cxbTm1/4kIDrbCn/H+pwHN
7a0s5YtGlSnL8OX2zHIPZeYfM5fomthm1dsAcJAcUjb2nH1twNc8XLywA06WcTtuD0dDzvsopYrD
HaT7vvIW9jQvUjtnLZbVmRvU2DF4wcVQtiiZhebfWPozou4LazQjK2n8W9gv3lWcBGiADjalPTdd
st5Uo5L/M/8IGrptHOYvEjppJnyw+unKilYEa07X4CUTBB75qzo68X4LQwJyw2larFfkSlD3gIQG
dDvz7144rQyLyRbaSayFkTIDcR2G3j/LSRWuHEdRcA3B6N2EGBmBpa/e6p9skSa5c9INg+4eizNc
5gIsCQfUrq7JaUJOFh2emloaqOE3GJih7Ay2mvwr1ptoguVankFs7hbt4j+icg0A0wbeoInx+Pet
87t3yUpYGAifUQ0HNS6saHB6VeNefdkJYJQDQHSFM3mRmdeTUwW/8Yz87MiuLlJO9G68RQcxByPU
7UCrWpVkOPVMjdje7WiieKgahlxa/IWSCS6M3flQWG5o3qsLbRYlVl6tYvXV0DbQDhJIvM/lRyz3
84tWclw6S8kiKAWdN5fTA7gcwctXh/yXrTwWIaUZDzW5Kw94LwRfExy2mg7WwcuUwLjlDDXJOrIU
nFOpjeN8C2qerTWn+1Pew9vtBSeO81oQyj+mgxPy2EdiUDNN7N3Vzg9qf2TxICGzbAqB9T48MshY
ybzf3k1ggUTKshNfppVF8CtHOtnty1ZJtKdrHTXi3I/B3QOCcnPEj4xF2vYCrwWOoD4TLclg3dih
bA3a5JRCuPd0QFdO7Cuzkuori9X/Uv1xnBNWzHX5bPMrPy/Aq0iUfiUVTrXTeLo8zOM8xMAwZPWa
hAMC998mzsPUsjOTtj4a/zBSDhJJ3AumRTk6wefWsz4xxwmC6WkOsamNoqjnopN2H+ghC48qyG1V
J+wTWm+2YGrS7JffmBeUChw4GLDBmpzyaoUYIZq7T7l0QcpoITvLCcMe32qZRvUzcKpriJNIyzR/
aoE7m0kMWaWQ8gOsy+G0HMx3r4SBaLvhC+7pG6HBrpix9yELvr7EiCW1Su7j4oe2Oiz2l4k0zXz6
lwuoXjP/NoO/yc8XHo0ESaDDE8peznNY0rGAeGXIyo70xbetL/GrimRd19+GDVgc6SD2rYWe96Ef
ufAQmT9cehFZQhRdud00QcKN2vwlMysMtRr8YEZJjC932OKzMTikN8Y8kHOBh5cltzaM4lspP0QM
Cfm7hzDt8THe2jU/EXBOcXxwBcSFgcyt2u2l0M1hwx2R7RzDe3UKxfeg2JFb1QSfJx66wlJ9Jjm9
S0cVB8lfWyesrR0VM6UDewkCNZ2I/m+4J8eh8eIERKYTO98FQdNl0KjWPji+txUaJ6kZ18K8pkqE
1v8WXxCc17fKIJu5qk7m4L5U0O1LTbQJ9rEx3IduuHFuMjvbsirb+xPH2auE8ACOpjd5nkn8ixVE
o1WBP+boaJ//2jZsumOtImeCXGffx2azmu4n4fZtZhhpPNJGeUH7sSmHR0p/DdmpN8oc8icnqrAq
NWrSGlrzbFmABJ85xMAb1ORXBLr4ouoj3AA1xuCr1Sce/mbd0ByLjk/ZtJhtItT78dPt6qRw8vo9
aVzJ7ayM6i1OzCj07VYHljYG6RFpE4kp3yiZn9l5zQC2JxKBqLeazBcgsfmwl47sp77aZDm1ECf9
Ow3z+hUQnPK/orgY4aPeYNmF+DRC9GOC2phOZ89EnqO+5JHGNdiAjUNYNzjSH5D+u1aPMlRxNhpK
aUvK+IREpvk/1eTRSZfLH831rM7Izge7KBn10Cpeec8aYZJP4cD9zi1g6CLiv/RFfZRHhOF8zBKD
rinCY3EeqLodNhGBe6H77tnJXfMXxIXmnq6yYLrDnOMqCpe91EjT0brGRglXlsJtBjH1YZSupqja
F4rHhIkoNHz6RhJ8zx27Jt7X7/bTsNd+3B4sqBZHexyG0xDO1x/I5fVIq5ttPSt+Z1r4OudfjK4D
Gkb7pqAt9XuY9pJb4C9Ufg8IsZbXmS9U1gKouzAehcgy/Mg7fe5GN+XP89xGYtU+6W74YhSx4JxS
qbBWLu8gXPZ5ZoS68obDpRaYreBrKr+okHrK2yE5rRdJFNRMRvwZvjnvs3BtNSgDtOBUDycjn22Y
Y/qNDfHow8aUoSEbLyQxXpC0s17yTHwJiYAswB04MBDmcNmjncdtPEHanqbTofa6jnmmjRtiLzrf
yJWM3QKS21if7+u3sYo/JlZo6ma2Ul7Nu950/nR6Chtkurx131SDaQyBTKFrP/XDzcmuTThlSqH9
xMJTfUd+ujidGrKlBHFA9TB74mmqNlPGH5rYBczogSzmgdk97+tBWm0J5SrtMVY9+NHGQZmfUvwp
aUO8gVulpgrAFyTMAVso8TQ4pHItawgMVC8xev4sphIPAfa/D5HIOBGKWsYtsrJCK8Rpxe+Gcs1A
2YI/G5sMD/4cEMlUPU5dOIv4T7ZarySwnTochS1TPW/WNmPT9fF+Vurexa8nkjNGOGcXlMH/pFyY
CynPWnQQwfHLW5BH+51OR60EXfzExe/rlWkYQefwx6nKBevTyQGlYVuAgNF/JsTeSgOCuzIaPKc7
6cxHv3S3CjINISs0nrz6db2mj64lkXF/vaCAsi8F3SxmhIs95oIigvx8d42Ullr6NrCYq7cJSECE
x6aRYVoDmIF1j/zkse6Qt6XvZYnncJUv0GfrdTKgOQ2l3/6IuMVD8yniQflWYNlFMH4meVXGxVzK
gXgOLDUQ6pHkZmZkFEB81S1wElbZqfRYcvRh1FmSTvNn0Cki1J5qcHORpkIHY5T3+QRrGEkPUUt6
j/nW0wqZh/1OvlMJ3tA9Ms3eYTbUE5g7oqialv/t7GsvBN6WJMrOs76pjrusqPIn4GXjTwapLY9T
QAspo0S7JcD3zvkw58fFIsdtAiKKgRMM1toqr3v0GnRgJxv2JpfmN7lthBoF5DQbj5YSz7V25DMc
a+GcNA5nIAo3AFHPgIlWUP28kk4MdEqZwaTW2j3hsOiPOrVd6x7Z/3zqIE6PZ4/+FkeKJMTBP+m/
ZUJ8fj7sen34ZU8Xly88uqV1oD85j5lkkel5YzRiXPnaHl/6ne1G/ToVIjU6im2bqGwuE6tudgRm
vF3F86gPshwG927aOMNYrZJq2Bn4wx61Mc3OVi6UkwWJmsnq34HsfGrWiAgRIQfxOF2A9iWgFpGu
MAQIrLtg+4lz3fSPQwzgk7Ac3g/PCN7eMVTRJILZHTZMP1S843ou+wgg6fr31goxqcDju2BXW6AD
VUT0HpXBFjho/adcYqq1WRG1OgdhA6wyHiyramyPo6tu5HIC8nccyHaDLBRNeRDBh1p8qLVKdshk
guE+AGDc5OzzVzXaryAJ2KVYQIq86FJHBEd2AOV7FjMyMjVvkWq3i+CPhop6NNXEseWY9/TrUvV2
YbTeg4xdbZKkY9RGeoaM0Tb+/ZtreSjP/5ATx61SKLcAH1BMrxC6WpsI0NRb+4C65kI9Y5wSbBcZ
7mmMSInI+lLWS6rV7P5ZnekwE8SXUZVowPXHm4feyteP8km89yDalwtQvThKH2IPmE7DC2ZPSkOg
MPcVBI0wWrwvuZQH3D/EehlmTub7+sQkjOIJO2O7566u0uBaw1HJtCUjHsgFhpStP9gYDwovjGM9
2XkkN44FUtODrN6BAILvrEjytGUBZROWYU1CK2QzqZYmMUyBp6/KB7sPzSRAaxYZdACOj6BN+TSE
JBhxJQcTxqy2aeEHETbjJaOeivzzoaQOmj5KZimqo1MehxQFcHlT2TvPQ+0cfhL1XZpUhXH5MrrE
NVsysFtfG9vWqLmsOCl/zakOUEs264nuCxtJ2DfafB0e2drOt/RgKypnbV78y0uEG3cq2lIoD1bT
7qWjKwgDthvLfLLUXHco8ao81vE13z769Wws1aphRPeKe877aGYGiZtswzfSWqLj/j0eAuSlz928
ZnObqjcyNDPK69MVJr34/KKfBw901BDzkd0myxXziIXk+rJUuATxqXjerb7n6+lPA4+7KMly7kZB
YAI7czu2NPMWgP3CFagGHuYZlwjGvd7RDSrAYoDgDw5n95NP4K1S4kZAq0230P8hpNQsuoznocQF
wJQ3TD/ltWSwJlZ06p1g8Wg1xoCIs8iaztSbTdhbR3DLq4gz/S6OEhoWjfuUHdHrx44joqOs11GW
Jt5tjqqPBxDKg1aoWlW+wLIT9VFB5V9+hUidTmjp++RQc5e9F+p53GgsTWmLWykkJ+nj09mjwENg
5fE0gvLAVz1dkppnb8b01jkat38ySevEUt7XOWgYLdp++VSoht8cg/GOq/uIxEBo5Mw11h0DrUBB
5Wt97qoTQ45d8iKTf5v+Td36Pe0Br8EvXlGG5LNqgMnEeC5eFKcIBsMbzhLl0JwY3xDeKdw3VZDv
cbolNnT2Y+reX/eVUfg3mNJsjv/EiqHizNjzhxfObwU9yTgGxC+1JsDmEhxpgmSv8tBinH32Ak7Y
6trc693phl3mWa4taloND1No7XuznbELvIVf6YhYdl02+8AEKB+0rKg/LlUW92hhEwIz/HpoLycv
MDLeq6gfxAsgSRiZwosHsp1yS6d/mXfm5P0U3kX4PMWtpU5M+SP6KwD8zwx58TD7o4mxrLeD1bOJ
xbC9fvqt8o5tcmyjigeY9xaZnuC7RDkGDauDSW16feCfSFZmbf21geBEa9vlP7xiTepTmhWTZKpK
nEXomcnHA1HmlT8Gz0qamKmyZL6oaviZ9hNTHtLij4vGkiR65EXbecQ3Ad4tQCw/tjuhfrlVijoR
JG5eLCnhye+/uqNhviwGHuS+n/bg7L+foG661vQISCZDlhgAuVYpJj4qj/NwR6sVnJf71sDCGnu9
M47d0AZ8wTWunMc/i33Ys79CGfeni7lAXHHmQ9qUNeszupGnPMluTC46Hes/gG7aBZSiDQDfhehQ
btd/PXddeFD9PfviD4RMfobO94FpRhdgRuTm+nkd0uAz4aIkJZ8VHXG7T63PAAYIUi8nRjKQGEh2
BFTxpOD5KSHpTd91WAvexw2ZqDvTSOJNLsTF0mRwpv19fTSYITaGO/YYnlYFIro6yClpvHlYl6E7
WXIId6+UrrD9GhkwZllqJodE1NYOJQ6C6Oap7i/USwc/KQzsTq+r2NdB7+z2wAAOHVHWQe3o4mu5
Oay4Eqcvq2KYEPmoGO4u5xx8wfKAQj9JIJswari6AnRMmKlxL66s9AVPZCnl6QnbfMPRC9Dem7zm
ehxIQxhfPbHWBc3ZDXH4IXU/E8MnZxuv5i7C008UEACGv+08mww9Vg2Y97T002zcVP6ImROWf5qp
2hS0a9fuxp5avjgLMbUqVOz9H/BsrDGWr0scOWwoxsOztzdM1BJ9d+wvzscRz2XupXLhUUG93DEK
SVfun1sX/pToPHe/mBltY98RvPQt//I54B4qWJMYV2gO4i/ruWsIuZPVx/oOW36bWWXt48v03PQr
TUJvUTUBaTYk5qu0QEOvyv0AZ9eCXvoSsx4lE7SVnFAbN2R0GkW7Ct2o6qcm/r5C4xPiJTRx198e
iG9XTxy12YE+JIyJTBvV5p7X+XVXxV6Yb/1nHHrzootx0WotfZAEARPkDl+76sDJnTdmQTfjIdu4
f9adCFL6GfHFR/zSLwDQdb7oWBSVOQmSBPIfmALgd6s53jVnAfSENf3UEm+qx07euoBBN5D55CXV
Iowcj777vye50yJ3P/6eU7AfmEV6Ox+g0O8hg0PIvz2YcHRG1LHfHNqdXg8NXgn6g3Y3e9QlLU+v
svgyf1oSBSvsGrEn+cQO2770qcToma+f589XWwyiXj1PMsD+h4+e7V1iVlukPXvJoGyMUIrhXP15
JC/ByLZw5y8oBZ6jMPuMyBt6j6fdPrW90ufrwMiC0ziubKrpGIyKJskW/6sLIsHjiaH1HSB9SQ3W
14N3FAjD02FyYp0bR9BcQ+wSyvwwm9VFjVFprLZSXRbcNbD5E1qnAU1cSNaoRd2QZwtOo4rJbgkm
Jtzy339XC9NAfq98U3+FlKWWJLx830Gfp2hpnKMi9YrYYk4gVPB2ZbFIxMc4y2w8DSnYC45n+gxt
8AJJTwuV8IB2nzpknOaqz95JQ8MJyLojvOn1DN5Ky6fDYvolVCucENncjcHe9hM0V4ou00TVXL8j
AP/+oa/+fw+YiOH80dqwHntnbE96eInGvQDjKkEhbR/CXg4LgkXHFH6IdB9M+B2H4gNu2Nvxxzok
xzGauxgwUQGyjA3gm1H8JKOsJBeIXsP+xCeoyK0URsg9pXnuiXwiGTAaSecAJkQjEgfbSyYeh80u
6G92eRkJQLZkRE+gPID7W6nD9YAJiwl2Bq6QIIVVbAoJeWysGzpSmqIvbeteQaNuObctbns5IsId
M4SicvB62+5MBN5DvMCb+z5aQuGN/hfiG4ggau/pJLlvINCCq0tNu7cEEcfmrs38Zupu7qz32xq6
MsjQKkqAZATPNHnSqVLI28+qdvvbFybxalsX2901c1sKb8/7qCfc6bicB9vx2MDJhzm4Cw+Zhek7
fwBdv7JBUA5gI1Ig4+U3R/2WVP9MUWvVHystiFppwOUVBe1DHDeg8EUza63d97TeDGu6y0v56QFp
Jh4w1i6sQybImkYM2xk03rujwdY375TDaW+2V3HsM6SNZyRrFgv0tI8yvP+/z5wWbwLHrMz9pNcj
Pho5O6s0iLDBId8e+Xsgmdk5QtDRbwuXQWUwGZfMPjL+iVkXMrfA332lIrcNGF86evsvuQQ1Sl5R
isuaGI+k5BS1+B/ObUvV7F9quA91TI3QFuWLrBN7j3IZaBnT4TXBKuWGwtkZfREUzxkgs0mbuGVw
tuSXZMC6qdx5WotqWxhmjo9jQVTKsVQp6bG+aip19PFOSNeAV16LvNcCGj2fOQJwDLudkrH/hTvN
SXPdTQYF50x7B1mvBzwkwLXDCcZmh1m7O4Oh+LSuUp3mUhSTlX/FbbvvltJ7wYVVOVfSgzZpVEc2
RF7oGSg8sB87ybBMOEkaiGNxijNihs1yblMf/gw/Obwb2lJ5fNfRP3CgDI0gXgqd78yMCPMqE6GH
vCRzMkubzwGAMTYbG+/xkfYnBm2MS6EcOepgYbcSZODMyWMdPBFw/m4cH9gzKW7FNUX1PeGWB4C1
EOfNt4ROckJ24pU0tw1cjgnOAkEMDSILsWTcUGHplnPJyW/EPyBC01UC4yX+yfHr6QGgpVZ4o9Nc
1N15FP0fAhyBhoFKrLCQOSrQ/FcaMa+y6pRg7mLRZOBE2fPPIE1ZtH9BPQNHz9iw76RqfF8j2+Pc
KF7pARodJAypAhLcCOYrvT8/RzeBjdtU+gXGxiQ33qIeklDiVISrPf3OKUfCGSVcniIqYQOcFEAs
9oxpaLWMxJQ1WDtWYDjTCJtrdrPOIfYkMURuUIBEO5ETVyo2ihEhXp0oOfZ+TqPINFsBPuuqk7/x
qq3IdTDlzSvmFSHWg83p5XmYbpH3pTDax99kN08gMn78GVDuetrwhz1Djmo4MsAIwQPcJLmIidSA
Ir4udgGGlJz5pdAc9maBKJJRIcV/Aep+YiWdQ7yBahtL1/BsZLLWsOyKGFZkgIpmGp613WW0ykCx
ZHQkXdsQw3XWiQGtVP/dCq3eo+ReqJSPgoq8YfyXOKOek3J6btrUzhSzl4LKbRBXE+agaPXFg93X
G5+QrCAGEy9uQNqQwzxu46UeBQfJuQeraptuzEk1PH8Nes/sgHxsz7wXqqPzZUfiaOewqYUet0LD
8ZztHUAWe1NYWpDu6tQuD7eDBGoWsqkwXCNv7kZRwZsdRFGMYWRjVQ9Tt4GVwzmMvdfi6XyRLAsl
j5Hv3qXdbsHJc6YuEgBqKOAjQmKoWR+xknpraqoKqcIJRJqZZuphsjIK+Eq4zaiMBTPzAMvUmk+s
zftRGGZt7Udx4e2RpoJyDYEBxcF235k2g4iGK6xaXQz/qAEd4E1tOTFzTSBsCGcdpyMsRbHkxBU6
xSCD5aZAIzR6bwb7fqNnckj0/ttFhwnh2kx3ikFnzaQ1qSrk7yeNgucvD3PFJfRGZsQoPLBvegYJ
Pghr6k/xyDxH9cG7eEnSpYCZkU0Inks4CxptAScqN4bm96wtrAQ2Dj/OXN8wzwkABcJ2Emmgy+lr
XPNEtw9lJPmrXZeA19KmAjF1bqS914HV0MkRQdLJc5YFu9mDtS3IiE7rRI0i0wUMJ0QfaAPu2Hj8
WkHIEve7dP3VBNWt7C6e+vaYynt8i+YMDW3jeQ2MRFGd/3uD5hHqCss3d4WdmZxuY4pZBMAmMXZM
BOVpjICxGO2NF/p9zpda1iUVjvvqdJmKJ0FzkC9E78qOC82HRbkuqPFKMlXVtzrrDAp7E2jB+smP
ydjb5N+lXensbcMIiKNTT30zztugE/fjfvIXgEcgUzprWnrNAwHI2m3JSihSGU/07NXOJqNPimiK
rIeYUvs0EwAoV6zlDqq4hkf1novY2+eKhfONt6Pk24YI7V6TOgvgpRnJusR/4JdkzRU+HuUkZaRI
QbZOFEI0y05vcrmyfuiVOhhufjfxdjb4ZLtLDnEQwjfwmBnYVkedx7OUSt4PPDrPc7f6eD0tnG8G
TLQ5ES5TQVK7GrvRIt4HDtJVVLx9gaPDQbyRxLY0CbbgShd8IdcsJDjA1GaY9YfvJ0pEJ/00coCi
1bdJjIGCQy0nXkvQLfMSfwV2YgK+dr0n9hIlG++VmUZ5H8yjAp6EY3DTkyyh9899bu49XBSQxsu1
9egS2JPi4ZZymtQg40jiJP9xESaV1kUg9G/HnqJba9EkzOjdvnCCbhdM1UmtbfaXmkqnNDFrRBwZ
gGuHjjldys3u0wRzFFYXrumvntFPUKG3aKgE/HII9HaBd7Obvv5y2lxHTdQ7GXBsfzLzDUEjMjjT
KIQqoxA5WgkuVmnN9XDNvzye4PAdpwenGv0lEEPzpAvyzxCG4CrlbyzSsvQaizqHQG7tO21nXa+f
CyAZWpX05ssNsEdQfJyUrYR3Imn45fAVQ4CJoNbCTQdVEsBcE0VlRshHUP/SIGAKxyTYTYs0991L
jUU2Z94TK274n19c7qPq89jdQ74AlXK4Z0ynvUYfOVHxsfPuCBzh74XqJ28p7y+X+RmlLRArMVpE
SJ0aD5yO4hJ+V4XvOwu7tFmjTBScnFdKYDp0utYnlWObs31l/j5UVU1xAoZtPjfzO119SNQE/J2B
1f0NOwSl6qsJ75BUkfLtcLp+2JoyUF1ixevc2ZOETguquw8PDb56Ox6nK4PpE0/4cWXHpEWWD1di
pmKELHPqmNmW7qKtgcoNxl7KskOWRLrrnBobHtlHNQwDju8dlbNk7EoCsoD9QpbldaQe83uo+7mf
xn/A6DrCV3Jzbw+c8QBLig3yjeq40QmZAWWXheyi0NzecP6lpwCihlys4kVXWQ28fy4XTdBjK+Og
lrvbI1rvOr4s7VDb1W7DNbW71rYITkmYoqZTKHB6xKPGC34X8Ylwsy4PZj9olzxectt1LGuUQ7c2
7yESTcxHxgH2v5p22NUZDM2FuxuewWbH8FfflVRi5uHuRuOhO7irhmicBSFxXTaRzCffPSfDjGMB
QGufHINugIGkLYJSI4Ox5huCZ7I6Ge4ZTyjMYQ9AFay8SKjnPK2OVkuJ5GpQ8D2B/Itt/sBGR05i
Lix4k299b8G6q44c2zqg54p+YVLHixSEZ6qw+FSx/wWnVqVFxcMGLvDyQ1aUElFE3IdVyBd5euni
0rB0n2JI2+XQIEtKpMC9gKdppXATTzpgOsCgRMKPiXHvMqAAXG+uze9cHaAwDT21+V6MP0FrdW4m
ADDMxfI82QIFypICTF7OnWJoBQPN2gw6KEc0qyQ4HMy+vMvVtxQVE5LC1bxxzfb83ad28qHSxLYK
RrDxFKhiAvE48itJIIhUl3xWGh74MBNMsVksS3iUz61d4030iXtZx9j3N/0ZwS4uReKJ+vW1DTax
ZXX1QaAvHuGx0T7+aT9rVTtg2eeHsgrkrwI5Hj4DaMIXO7K2lmH89xo7fI9hrldESCjzBg5VtWER
6zUg9ek92c6LdT+8xEhdNZUu8y12vgx0i/pSb4lmqN0zIlQmwiOOvrprl8xl/Th3hi+qE/KJBLGc
FTM+FdCBPJisVxikwRxuDren9Lvf1KkeGZXn4AHg5kOv97OkAZKdY9oTbEhMuNl9FF8mliriGRu/
XIVbic6uFg3tN8ZnZsi90LRX/bRf3oJJcXUMK+NSiIaE1GQZJppN8kjpl/iOU/j6lZTUUNXRzek7
s7kc5/8QMQm/tzqUoGuJTXiWhFis076wulFom+prTmcYoHq2tBYzABz2s3Vr8qvFOy8lNO/PmhC+
MB5xosYquOMw1OBE+x2gGIa11Mpo2oQNdBbpQewF9/wp3EvFIyc1Txj75Qyo/UTluF5bg/OmCtCb
bXzKxObBCYDnzPQCKuwp3KatMyJlKN1Q09yY5qEY2n7OtCgZqGY1ALmUL6ILaWJGuWQqLDbvwHA1
GwSWLVnCP2EboO/0hY2gJ83dh+leB/dpXDYJPVq1DBx7nxKx+WJ2NIPqSWlnVsyS7ikupomm4kBn
gIEvcq1DoOZPkN3udNERjRHIEp2t85OiHJc1SMP0/BSTqWfaLqvrusal9B1sGZ4r0k/cgcqIF9Jh
PGk6iBZoAXGdEjgIf9xJ/hdfFo7qRltkqPfaMjMtPbz+HxeM2vINhApU5JoR/xHj4PWDaOodKy2j
g+T6FWx+qwucKJZ9b95ztNJs1THqBXcFYeXzpIxfdwA4vGJZS4Dn0SbY0Ba+mqqLWZMrD6Niu3ac
56Y1md6ZhOJh3CP4ibohpItA7vA0nnkz1fnDDeT1sjmwj6Nu7w5sSh+R4S9lQAxmswFfLY6l5u8z
UFtEAiY6dfb6qnHg1PQZy418+/rRhmgNeLC9vE87aZpR0xwz/FiQsqQhzrnzSTUPmQaQTXmvvcN+
0b8lw/leus1hqvAKQxx6Wc8abhIfx/HNpfBwiRGYruZoNK460mizEkvUOJqjAwjoIC6jRUt4xTf7
9WU51fFwBsrsgA73qZsSw605yyOVxGV7rjZwtpe+mNUubavK/DzpaRLNoAK2SFmqHfXWaoTwmnG0
y4J5Gy/ATXacE7BdLqhk1Cb1TCA1Y/FBecLsBBnA02hcECpD/veUpLhGpPxeCvQhgNvlHrqha5tF
olnHNhvnpjhDe9NfhOnlj3JxsM5HLGcmra33C3wsVJmac/oGb5MlgzxpekkyPvyjpYv6y194lp7x
Elsbo6OzF3/pzh+FmYKDIjRxrxDdoI3RXGSFL3xUWQXLJAqo7FCwMu4jQBeXCWD8/HoY+Sj2+MEy
BlaEaHa/EUlJ4zbQjT457i5RNdwNu2RsnrzCIUscq/oGNk/AE9tk+nxqACyGkNvsEKJpP8OTqkb1
Nm9iMEzRZSpNb+rO6S21uJnTlVG+pkJMrvqrKT688c+ICk92vr39oiRXuIG2RBBFQAfZWXYJexAS
hRy8n5zhIpFplB9NYBLa9nc6RXvfXqrfb826qjBbk4PBz8M/Saw1VSgLJWFyDt3aHAm0x0GqyIlr
OTQINJhybPxoOlMXkd88f2OyPCAxhhRuo6QroAPO+Echn1p6nP+bmQErevbh5IW2PcZto+tGJOML
FuOOHhi7UaM6ScPKyfSD2PR6di/MG/WVa7uaGiDAMnfu4QC02Hcx+3BRVS5fh787bvzr76dgEDPo
7ZX+F9YpvlwCxsy1V4Fp314MTkWAHKAnYgODli4LtZrD91Ii5kSeUUY7tpqIucTsVtbEKwC0bRSi
E6vqHmy7T4C0Sg2hA4JAQ/ocgqDLAgSds7HVPONgHHB4c1az2w73DWR8U++egmWn5kT12xscmk5Y
NSji6N7mjheC5Pbh5iRi+dgkNpRUYM/XGWTSHfmmcY+enoRnEyzRrjyfIYzp3tHFCUZUoN1b+IbP
LfAQWameuX3u8wvVKLBBK8ONiWSONAmwk/yVcqq4uDJdZMCYTw7FZ6OhiIxusob8nGUAqxYGfdPw
zlSEVa2l+qwa9j0GC5GO9CLEf71+KP7zW1HTCV9/WUNqPVkFmW0ApHXYbslUf08vskjMq4Cn02yb
7IdTI9trHQEnDj5WLVqkn2Ii1werFF15mIb09y75ylcR/yQdw5+91gpjfYFJox39R+JMMO06s3Xq
MH8+2OGXxwhRAf19OhqmkUGPimt38JxdqXN+FGjdcmSUHgy4u358BtOKYk88UsOEfaIr5Eafl2u5
EJ4paZsMrg5/+z++wzBJov3ciVgAI5is/BFrFAqPW1wE55e/vm9MUzaxYk6GjKuCyf5eaQUlNO5T
8G2olh7RlawvFLSeWkmiBDbcykMrV+IGv+1IlwDsP3ZKi+EVGT+C+8//rNJELxFI5AEoH4C5a0gi
Zle7VhlRUoLLGU71HBLuzovw+fywPcj0IjZqLHDohcVljvJ70ouiMvSzL197jwhkZHMuPU1/VQ+m
iYqhBrT2+hKW0JEish68fAkssN9hz9BYNYHaVOOVkWidOpw9ITlFb0JA7bxhaqmhc9tp76YZ62xQ
fSZmo3evTEbkCxPnFzZqJ3r5PzBU37wbBYADIHNCBuFi74Jd6E+nBc7VOyK86l0KyfEY7UO+O/Pn
RAyWhbjBvw6vcYtkB4um0GM7TCd1eog0bMEL52178rjcjFA3kZkUV9t6KqgJodd26k38e0BfLKgB
Ecc27wnUIzU1HEv50A5FncgJR0M0e85bCRmWdZ45iggpwWkR/KCuMaT8QeSlDxjjnqooGvViXdTL
h8Fja56ge6wQPyWb3hkLlRN7iOaB4ogAD6kBsJaxXEujPN2nsAWKQuQmje8NhyyvpozLRvk9ikm+
zS8ew7z48sAu/RaBW3OG7j96yHK+XsCnJAiWdk9CUNCUocykTU1Jom8iyIRcETcJpVcxXggxqQlh
JiGCH6TFlPd9sOpU2smP1MQGJcyyqI9aFnFB5Xng8+Y46fAi4szsHc/tr9aIsRnS7DrVe7hmwwiw
g7PpTgQ/88Yw5DGhqI0Jjg/qrI6KBGK750cLqBO+e4hcxjmkGOZNqpNW8yCfVtXW+t0YKluV5c1R
TfUm68ldA4fnS+tSNvnJP/YqwThpbXkr2SI0Y6W6hnDdKY/2KhwCDKTZgFp296HmGeL0Lv3uXJQe
WbG/t+h2icGeRrhCeZjdq4T6GZCcuhOA6fcRoYHUo57pkYDbuOkIzCtn7zzqEl4c87lZDbXECkXi
vFOPmz48iST7FuRAt/wJwo3uS+7cbeMSW+Qb0qfM0exfJmkLCHfB2Iaq5864as1wXci2x+KU4wUM
PWSbRlMzfP5cdRjhRLKxfIWXlbNgWzENzGj9ec92AGL5cVqXqncVaFes4WUrAixJeXU39LCChVjD
0HMYXx4znueVNrnWzAF5+bKWUDt28cFNoZ7r8PbTGvtMrn01/gREwXAxw0Q5aXRr80r4xf31h6Vl
nm8+gTNhvZQ+xTy2WiFm8ZW2F3j8cc6iUBaSmAuFceHaKJ4/gHnq/SepRni9sbzyepCFulrSy5g3
uKDaHeDBFH96P/uMtXzi0uddoaXdrUNnP6Z+p9RcQVTF0htSyAiit2aUpOFIZr3aldzzr09/QWg9
ZEDJtkPMDdfCQuq3SldcqIAyLN3ublGGCjHBdLMQRr2ROZdyrh/M+zMUtdRP6ItMlj0x2yQfLKY2
DN3PgNyk8egLvXxyUVxiToa5evUlX/FpJp0wFaEMuXRGZqfcJgazh2IYzhALFriHKKNj/lkxgKO2
kxdjwfY4g7YuGTDl/PLhE2V8MvOkAtgzoley9M3iQHbSI424sue0ASUFApYzTlZPFId4CiYyXdoI
vuAcqvzulZSIgpKmCzST5qa0R+nrK8QvTn0eWMMa7gKDgJLUPqCojMYzFY6kAM8zwCQc2CD+EDHV
e4/94jZx/OzKxexEjLq4zEwVdqVWr9DSXmift3DrewcGFhVggN1olmHEhK46DwzEbQFoaJIygMmX
JOP1MnVQfEDtXSH4pLt5gZfOp/Yf+EGITMwFLJEp+KHLTuM3OeBrtYS3k8KrcWiUkx2zpj9m2aQY
Pvpo/3Vl9hLB4jDQG9QbJiNfHjMYehNCuZtOnU1iC6HcDqV6K3C8jBVYRF6F5K4t29couW3xtKJh
BHocptjyUj1DEeBYaCbWFyor9G9NrDdTKNOP/lacC5FKaxTrb0SK0+u2XpDQ4+IXRaKJftQ6wXsv
1hS6g57yVClJExG9LnViPpLz9UaBksyHEBm+YJPz9xB47aq6N01mX/cwYw0YxMEcZtcs1YKtxZgR
rQiR2BfGJhVWSkoJV/yNqwJc4owtZYnzdSzmxe0x0M2tKQDpXMq42ukgLFTsdIxhDT/za/wbn4H6
WPiLhsuHSi+RW/eqlTrpHADQVtDzvi/RflJLQlgbF82QLvLwL9PORj0Z9GbVoqQnjInoZIFpKuQd
suNKVXZBS29DZf1bKB13mDH610H02/rfeConY4ZTb5lIPSLDDk0AM1JXhYnG90Uy7gHj0+7FpCoU
L4HFIg7ktbm2fW0NRuzvUxKPwV7iKvGne3qG/AraREEnm+AXXafSD+LeppEvXG4WCP0tZq3JGkyb
wBY+kV1CcyyDO5DaXhQu3gRNxn1cXIr2RHu5hgLzviLvnZnrDWOmv5Q6BPf3P/17WiMwLC+j0eg0
8gzv1qITUIQfNPzkEgMk3dJQwEYPAjop9HguTSk/3D5Q8Pdotc4Vm7BR6gY1TDfyISeP98Q26veg
gxJiPLv5i1MiHQj5e39/Omau04upWGODutMLMQKMAi1GoskShzXbo8zCwK7QKhAs2dY3CLoIYqPX
bNLyOC8fKffRzMKtx2x3rBQVoPSa+3B2Do5feSATI5ojOOsTBCd+9fWPRSKTU/2cAITWyQl6lGXs
TSsX5w69onz6jLJZA4shoizYF2fhCHvg2TOMRuTO8gHoNCknX6fRHFcE50z9sNcuU+gJoYX07jTb
gKka5dU0vjwrsRtoJB9otD1A96rWuPzq2P8kFvKOf9euV38IlwaK0nwtqrIja0fJVgCOfeC+/Yo1
edSv1PuQQEIfINUckzWhhq3vTIHMx36K8ot4CsFumuYZBNeH17zqh6R6bIOfAfc2T4Wftu01Aolo
kqR97vkakBJHOA+3Ymmd1fhn54zMR2I/qGwqX4mcpPLHnKxM7nXBfW84+SBETO6sSSRDC7lc6c5O
qnRr0twk5JCyfOX4Qt8pUh9AH3V3PdWxWGgXvABYEwXnKlgPM0xkajivhInU+Q9odZJbyW/5y2m7
+75SZxuB+TkGYXcpHTarvh8ioMjXTxax/4hiJpFBoD1k+Jrwz/QY45vLODN8OHQHsmnl8y7Tg1AG
gdRxPFxBFtxB97lrgYsEdDe0nMwZuJAf3celAPRPdxJtEEEYQqd4wXh7wswTC76XPcsOYIG9qkAJ
zGcBdPMzxTyAou8CoGcbGYHstGck8Az+L8Pxrh/qpRo9ZCfn1eWzmeEmXefodFMjf9zOTvKSQZZv
AEIKClObq5fCyQDI9POBS9EK447onVEd5PDlGzKN/aEV+XIyBSWth530oAQaZK7kIo8Z1jDR4MF+
x9tFs627fzGYKejBMrCkKDpQhJDaTK3k5kD2378YuyWUpq7Z4Y/KAXGjzeZQB/aS2+h1N7KKQazi
FF8HmL00nnA7S9egaytp++lgMe1y05EPvd1WwHX2vTgfCvHSbgMAKIAks6Gw4ynW5OrYNJylCtsh
MHzrNDyE6znEeThuDqjFIcyZV4OZMa7W/XLty7rH8iCkTAaJgS2GUlR9KQxoh0S4gWRqteCrPU3a
gVQ1wwbB3x51d03LEK2w+GzzjojPF49PvqS4nlIxDzymt77WDz3teipeBVaSTAcMxvG1ni9v8cPB
O4Js4D4x9+Qc8SGzBVVg9KqA0nXAFUN/VdZISWVBRWDdIt32SI9PCELJU6T9H7zcAQQaHqHkn4Ds
i3kVH6l4TdvGwWUNKNiCuE1Mdw1rbE0/MBOZl+M0coY2FdtNABuAimPcTz228D3jHwc/dMCDdPxa
ReO/Tf2fXepXK1inGxdgy9YOobiwELKuR+0LIFwJQRxWyg7ljDwOYoBwreuub8zjRqzi924M/iIv
nC1uFYqJZbzdFUoWgllm2LgCBU65r0TSfhrOMCDXdF70Ge33E+IJyoTRg9Su0FOoG9fi6NpjuNCl
mdKRDcoPcp51lfl3LnAVDR/E4O6UGLez73VGe5N2nE16TfBDdU0F6Oc1Kpig4gk5ClYxqwir2SK1
Msi+YeZHX7ui39ftzFaa0BV9qvHWRrHKd62T3OmQHQOKjRXXrH7MGKz+h4OLQpuXiBs5o90iixMW
EZOQPxBYtcLiwQ1c/xjHbjr5j/w2aeD+gDyIvq+XOEBP3o3jOMeYc0LtZUFs/QNZ75AaZV3k1miF
p62NVXfC7KumLjwoAMh+CgfkdXCq9/Rc5AN68TAmSxfHDdeOCItpxbpkZbGJCgHsFR5x5NpmxcFp
JR/p5lR+2TjQGTvF347Qg7tse1FiJyvLH0XJiDA6foSgR7MPqu5+8mENNXKDJPto2eWGFBoqPr/4
MovwMt5DOIdIbrRYXFwHB3mCD1LfSK2+Qy+C+WYY/VVJvsFkyXNvojswLoQ1ynv8D8FNlV2nIH6H
wAlc/Q1WC3yUnePvvxy6mE99wBVSkWvKLBiWCZ+Dhju7YAZKQOsyLjRNCTyTE80+wajkLweXsNpG
touMhL398XmaFI0v3F+1b61zyTL9HcAtwdzZdmFs5zK6NLhEtm1G0TqQ82S7tx1oHvsvjGD9sjEw
Bhf7xRAkuh1M+gRXdwdkUlsNfPj0uplWQPq4Voy61o3BOvzM0+DwtE2yWKq1+zxXIH0CECpS6GdZ
OEVz6lxZoyvSr5sD9J6Vy6wMpfmR2iBUrgMoXhI5AAL/ITy5s+pGyhrOR9H96qzXGWmaKLvOPuiy
J0cw7IwRhngsXyFiIm0yIjN5dNg97Rm/Kn0F89jS4np0QQbVyBggfwYDcpaTPelQLhSZ5b5xVwXH
r7DtY44XDoWlHu//8TniJ55QR9Dk18TdwHLt3h7I6ZGsLNA5QfAOclrqdS4dr4MZJjMqjR6W+yTD
BHv48YYS7gtetAx7xVWYrpgThuHsrS9jaTqfNHrjsRbTLea9UOI6zDprjzOZcadnIfl6k0wQN0s+
Y0JeGu90wBQm2NvxX8T2OiJhpCWL2MNOdxKjluAcjlKfSDlnj40RvH7HgWHLM1x9jM7y1K+d4c/1
67sImTp52YGPEVqOwUN9yK6KQVKPAE0UBXV5cJ+zlLbwgiA7pYHG2U2muD9xFw15ZXfcb4fZlhL2
V9NLr8OzKSCvgaA/YiOwz0F1tNo0/fkZWBxfUTqOkLdrC4kN6TdEYzzvUZs7zO+NjZDvStNI+u+O
+3BNbtHxVXOS77XyE+sSrJHoWtXJLcNUUTyusSw4NU2TG+qdRxp+A0113+GfZLxsYYsmdpN4HmkC
gxoYNklPIAvuleR7ievuHhjLfCTqGN7m4jR4Bj9QVEyXrSLmlHT7cP1GE/dxFs670oNk6TK+U1Ow
bHcY2JqND1zZ+hGC0H6OJK/vKzdCUs86CkxNnRHI5NH5abInXDadRjt5MGJORM2i/15kB0xQS45X
nbldBKOrVNRLDO+Cuq36gKdf1zkJIsQ4hlxQY1NxIkFU6FO1DXtY8f9E2HhuX4sYjJ3G0eJJZicf
xCxlDG4bA7dAByVbaDH+cE26wnMs5dMmZ5MGUjY3qwZ0D/K8/PyRd4XcoT6F/Mgfu5pI6ysODqKQ
Lnv7sytlZI3GGpuLcFEJ7exz76KiHSESgg+KxMH45xe5it1piQw9efYRbYblCIAGE/VgvEP9WjE6
iVWhnrx69fdTz7ijwHRC+38mBiSeoyQJ1FL1piiL4TqQByOH2qrQ0c8wp8+Abp4rXjL0zc/SNuRk
Fu+V0WoLFrnj5tjKs61W4RXVHlwmjfFK5kHFPlY1iMFe3me+Ae6dh4HsZ3cX3v91RFqCvQ4P8I6C
tWYXeXWHsl+kZeN3cvazdFUJ4ioqpMWdl6mzBYI4/uzwPgGNz2K0fvQtXiBVbHDsB3pp+PbK2j1u
f5eNiO/PgFALiV0NA6Y4QZFp3cUuzCM4AYJZzuA649j3Xl3sEU9r6Zyp+R1RiEQ8PLF7fmnNKmtR
eX9YtQaKMg+0F6V5PpL2bpEkSOMKEr6xGmqzM32qTmb758NLcd1/uxbesTnkCE/ZBSWWS+XmJjAS
pGuVoQJLb/Yyu3z24cujijIqeRZtBUipe8t0eVDPips56ITneGVKCqaLEFEO3ypEN48jsNFgDv6G
lCruN6C3dmUXl10Mp8CKVMRNVTfg69Uywm1KWRuRYFT+gxgWg96/3WO6SU5aKe046vd3mqil+j0P
a9D1EnCQZ/E/2wCRZSFVn59bbZraHVNzyrKmbGzD9+nvpqZMdXFbfhQGmiUw2uPBj+FCk4CogVYN
vXB3ivuIuHw8iodXRNgEXXYWR3RZKPSlVUqeID+MXUBIj2fHLuUH7GP2HFoHDtolDycW+uF2Mcrr
cjPAHqqprWZsuNuFSzdOpaSZj35fOaVKXjucp0X79LGfjrF86UDdWhGkoITkLPh47KKW7j8vJEjP
7RCC6h4+f8QOrmgO/K90oYHPXj7f9CRvg2EnB2EE9qBa1b80CvJQI5tuDeY8LsZldCgwvsto+08b
sFMopUAY5uDNIuoyzN5QkbSeYesjc637Rdlt7qhds76KnWLrC9EYKEXRM3fpRPpwrtZxoHOCjb/b
Ek1C6Vb4E8hWt42qZ4chQXzAw5c4d91Fi4t7LusH1g6XmaHdsgfNHd6u/ETBPxEict8uKBYCmciR
0LsVc874R/j+NaaOIvenmhcUkMIJeVtDquan3FcEWFuaa9pZ4z/27rJLmy19yNs479P9kU0BOjG0
NpjdyZLhcBf+/jBLP8w7nVcspSSKK4zWgiZOwhYsF3RzSjMvTbc9Nl5EkMJ249SkQbKDKR7YxLsp
ISqps+tM1rvrKMVWxAnYScOGHmhzInnvalQfAmeN5KcRn+tfI2y0uzK8x2+tUkH+vp77XfTG9Bxa
HHjZskj/6QVboi8Fi3w5eP/7UIIQioHkbX+EUhMDZvdXS8LJt1gvAIgFnzSvtSX26JlcmbRjuuWD
MXF0gERSexBvhKt4LuSOiIz3f+Xi01CaDpmhqjRmcNbQs/X3Cxmv0FTQoSAzWCK1SohrZJSpeM92
E+cQv41THHXqBPz11PM8EuExCjjpvmIlecwMEoE+PiLr+I2rUUusvWMrO818I/MoKIuigzzDiyZW
Lj8Z1i4vOYe4ELtaZK8N3eldrTUwZypt5j321uPbgeIZys4rwlp8N0RqDStyEqL7po5uW/U3LlDS
UTqCUKdumZ8WIoNdyj27cp6VUMYDyEISoI5xWUtHNgdOmjnK0gv9HzaRrWx/CJZ5rJFiccSCkmfY
fEjAXSlT1CR5+/57LXgvVp7zhO792r+ssm6PQYfo/V/06DOTgybSvYAe8qrODGCHg9TKuKxELBG5
xwbYTyz3/+LgdE+/w/GYfE7+j9yhsHEMW7/6hnLfu/H2+yMrkE0D2NdBv4LmKEB2RdwfwqldxL5D
Qh20o95yiShMhA27yXvgXEEGEbP+6EYLIkof260pm3Q0mA7pXtG/Vwxr5nwXun+EaCPIouA6JPSh
JwuEaCf01ljNVcP9yB6yH/cYQw4Rh4rbolxBxj5fTQ9yBDS0r973FSl0dAYhH+jpcGA5U+iidjU1
g9dElIdYknYhxHfSgRB2SVGFt6wWQKABBiiZunEVz1i47gDJZre9xf7W7jEWHFvm1SC7q2xX4cLq
jqBc5GF6Fl9jxQIeCFQJy89u1DKT8mz7YDRgTK0zGRk3OuX6ZC5HS8zmDWZK2e4H2iiKQlfVqx8Q
Bhv/9mcieHfkZ4I6zvmmtzyMgdT9yXg8FnWL5jRmA5MfsP5c0RlD6ywnkRb7FOp5MqQc9gcpx9SN
5ewORYa8OlbvvshtjENe6pF5jU+oLMs4D0TXNeKGmsz04Yu4hu98G8fWohK5d6TAvKGP0RgH4rLf
lGIGT1yQLl48e9nYTVBzzhC0mx0gwicr/wh+NvIJ04lnRVJKJO8RxLZVTVm1FhLFPN393fnG8zyP
5Y0/aoWT8sR0TEO0dUhm1/dHqd5qodReuR5uVRSKntsDi70ht5AnWht5Za4isoSPBgaQUX/Y+nuj
HbqBaQaaU7UTl9C81SPQqTNveItFRGd0lFvSx4PH7uNtGIRtrQC6tyvz7GLixM29KtPlb0NeqH+1
C9+kVBtv7ZikE+37iGGBTSRElDDm20VM/ZkCBZiBBL8ujqmTxgTczn4tsz8T15tdlhLOcVGfBd4F
Qyor4TkI0TgMJkirb0S4fP9EpUZb1CaAFIa28Pb5uldZnnlR9keJTNBeUIsQIqOnEDGHf5xCdGCl
GEb7C4gErV+GdtCOiaxLBCMqIfjtpMChAP2gxaztq/6DUtPSEenea/o1Gz30nEWoRlRM27dcBMB9
IulKg6QggxG26RH6JtriJgNtyQBE+SVkaRH5wGpcQQepVZ9EJQX+gSci8unvVemMCmAsf7ZjP+8G
FkJcDkXX70znz5maFAvDeQ3bH6OGk60PS1KBq/yYNeNmYHHLuJd1N+0rvMei59QuIUzeCDbZr9mo
ro/W/X9APr13kPe6rW9H7qEFi9IXoqrglMso8ptL3TmzKSlgl4Di0DoCuPIFcHD929+FBzVzRIK2
8FHA5VTbu7q17YGNsQ+JRcfcDPZngVAmSMqvHnqagoOlKwpDZlBh3PJNspzfzKXchamWa4REryk1
j9vdeOLFxVd6zQXXVrCC/kV6e3BQz7DLzF9q2jgqQ6RCR0+VDEj4HcDdDaHDP4Aqw3cwEW+F2kQ/
NMgyJEY2c1lvck91nLdWl5h+/AC1iLw2g+E02y1fjA3d3bR53HxwKgG+aCftlBQGrKUD3Hp9xekS
9TKQoBpNv3f12nK3deO3SIUh0+q5nO0wuddTgve39I/QnDic3iUHsYaaATinGAEUZUn1LzDIm9Gf
XRQHdoGUIRsgrNnwHzn4ANSabapzywpzGJ5tH/B/wsGSmsqMt8D4HUhZck4NIweaRJFSygz5HJu6
8PoNpCouHoaWrM6nJLltQKcikBZXknMHJA4GdOwkOFykTjElj+lel82q7yw8UF6P+l5UGlD5Y83V
IanOHnFD83/norQ2FB3i+IGhaDot/kEO/Q0te/mEO2BBGa0PzfJZx1mjPM+JOnBp9j8NCO8BfikL
KCGEtwqnY4Srmt9Pl98AdXk37Gwy6M636H2R3YM5Gi5bkwvMA+wXO64lJB/YYFGMrp9ICblbiRrm
RDgUrgBLWIGG8efQieKxjbmvb2mIjt//k9pnx5RwXQ8rWcvLACXEtMAu1J7G8B3Yk2DvwHeQm4Gr
m8A02osVp3M7rr/DsMrYTcf/IvD3+V6wBNIjsaIXz82yWS7enWfAeQFqX3P1a0WiJhvdIdxjG7kA
uWPRbZ9sh2pidG7gs4SCtx/4xCpsup2lmIlp1B5IaM5VI90TfOKABsB74/BkF2V8hh+UkHt3ibc4
eNS7TGzA3/vDxuUTmNV2TzPGMamttAjizyCz1TIPNKY89N5aADxLQATy6Jyh73wG51JtnyysVk3m
yfWzDgATozx0/hOdutzKqQ9A6QewI8CU0w8LLSMBWIS/g5IM65JX8S9TMTs1l1jYkMLUc2L9vhNY
lfY72wlnsMIahbkVXboPE7HX2Sgrx/cgJcMjDnZkJ2SwPZohK9afBGmAoGTIzyJN6lcLt5Arsv3m
UJs9R4UTAJUHExMbCO4jaZqM4/mBFFoZNT8vVdfbdy/h74GYnmfMOYGlH9VRG27izdNrsDucu4nd
aCHhmI/NCN87hGJxhTfXXigwP1RGpBUFTnxokeD6IV2H2OzMJSh95rgOZKbPJX536OTYdHaRF5g+
n9tVu3jG2Ylkd3R5ITLQLeOgHVjnTKdPMWkMGfBeIuuCy6PMZ9y/OWjYAMTkk+mUVKFzNwzJz28W
sDRfChX6J/JP8sKSQ9O2oDvGwvIVmfTSLPY0Ky14GA04wBDoUTn1HcMfCZvzhSLhANssTxoi43vG
JusO3G2AB/ub6uJDOgohBb+svejGD2kiSovK7bSdyh83qVl9Bd9P3idUhi8TTnopzOQxwuhzT29r
5iEdehznc8RvG93dIFdfsWtMGBUomtqx2w27C3t1o2TOrNwdCZH0mgdJb20OyB4ipzE2KtYB3lbc
A7vKnDdeMzS2kffC0286Ch44BLmK1LgyiF7UMyJn9H4q6TCuCc+K4jbRR0oV1peLM+Q4A5R1blXO
Ih1/rudQdhkLqdLnDsiBLhm/Utwhsc1oA2qC/Scf3alkTEfKGzBV9dWe7afHOmalyyFM7Qm1MjQI
5nWjHGNHIzDZqA3LSSeI++IreqZdtjKj806bNbDPFycLpOT5hRf/sgvUvyDN/8pQ7q66TS/rDZRH
eVoHEOXVTQAhOl0zMNIH81xKLgPHt8XnScKTdfXniFNxp7y574wHTIUuMtucIP2zMN3S9ZSYXQ3F
v/sPoF+mO8CDqASAesNV4SalC0ex2E1SRd0k2DWeA1L8hoT2E3+CthIKeQ2994XGiiM0zOgssDhO
QjLk8W4mG/wFH6xh1RcU/OV0XOz0sqSEcXpFt7f6ITc2uiWqjgbeQhCNUzxDECyB1of1ceR/8NKT
IKwWDUdfZwEwibJvAUqD4Ua5WaVb9twe9g/tpscqgzFVMBAg7fJBe/mzlzsPCi9asFirVcsg3a8G
Pt7UvCwQ8JbH1PLUoxvryvlyO2ra7k4cfkM3TpFa5YK4WGiY2ajIRPeOybqT6ovIhYv4dCYvCMQW
+54JjKJQa8bCcOQXDm33Y1yfU9J3S2MrjTFWRRq1SVuRqia/Xqx0wRZ7ms/Ys0nwscWQ7qBkobw/
uzSTLQmMbxQ45MNalaM9EERVx8qdhvjHrmaRnS4F2p+ajvSYZTDUHXu0vacCy7BQb4WlIzj9srER
TqD4LTpcYs6TngNsD9u5pcUfr8337SI6VlEIuXKr0hASHxQOcs3mHtjqAH8eRO8Eld2Kv+x7epF+
pNHUkon68xiSMBa9fFqdg226t/KF21r1PpMwS5xSiFB7C2PvmEmpdqpoyDtJnpc9uu4SA5ECOWBD
2oVoVDEQ+ZphFynsgUFgHoq1KrnYoJCsGuk4YwsyArVknGOh7FKbgPDPRlqEAo7ZDIUv/K+0xOjy
YRnFzDZ/PpUuN4yIDBUuicRMZl/92GpIeideIxNwu1klkhl/E9k8owhT9Rv9aRadAlYjD5b3bPVI
gmWVUExR+qxgwFaWfrRMjWmwCcTCNWCnaHIpfElQweOqmQMAhVw/DdfYbzBGPoSkgNYtoqzd6CiY
mMQF7aqZDGKzlSUdVXbjwn20UqZow+mVy75vRHuloXxz4gA9gsr5aaG8aaDBQ4BIWuCbWj1I6wLU
dz0nca/Q8cUYhsaXLuUqzL5OxKFkqvpGloMeeT8bOHrDveInns0mAH9RcM9rlwOPtW0b49DfQfdP
4+9/Q+F5pGNaH4mYL8NA5yY/qGgAuxQYanqITdCOtzEwyQpPcP2Vnh9i5bI1o34NXfDYQmEwADnN
Y0gnT6eeNqnZ8kR6lbxJvWipx/J3zO18EgeLAYJIQLcJGySxRqftnB9zLN6taKvZqUgTyPp+uarx
Rsg1p6X2/Is7olKVPooCQTXaRaKyKDOx27Aa3piCR0c2VZmlnMIL2PXgIkRqx0BccflHtKC+EhA6
I1vgmBy3tafYSEw4kMO3nnbIXC3PwBAoWIJF3u1mFgqAVR0+J3FADAxwfD5hgh0A1SU/qUIlQdnR
mDPjIRDvV0kpZCunCPsKZY9ljJCNA/7LWwWRMRlHckcklTaaWFscBg5FGJeMHEN02qL5MTlP+LPO
IHZc0ufcvNuwkP3nZ2PM4c0cQ1y/5qoRAanEVhDY07cutAXQrmoobcNqgVoD1n2VRuE2itfRcwKz
+mMlxw3bWV6omShxDUykDOlO/gGzsAdcSdXqZrh2186DLMpBgnCSqxTmgpQw3jCRhP1g8CXQ4SnO
sQyT8LPkhMruvRBoKUZckMfZzAKq+K7K5B/nZUV1Gju9i3EZkqKLEKtWH7g8DFG0r9JUcx8vN3AR
Ti/JWdKmNaloxCm0JAUmeL9gIAnzM4ssVtHkCwqg00R5UvAEsiuW1ity+HWQ9ATDW3fwYOF9dThU
pMDz7zIvmKmYfU8EW5ZIXBzL1BZu9TS2PRCB57bowfAH9gTFWqzA/HfIaY/9e30hb3QupNqYRPfQ
Bw/+uZLcSWhE3R/y+7gqgOXMD7OsFpYo/DxPnJgu/1yUvinqvjLCMDNSgnNNn1DDggfPQbIdxtDg
jZmubfWiW2CyFV7vosSbHVrNCdc0YhuhaTgL3xNnaNbKXBRvZmjpP+rlSQtcb5jaiDQ0gUXRvYOF
SGn6z2XEKvI976Jh0k6fWVGvWh3LbixEQnNUCEXPviYqziGWKBgXZQDPTxdNO0y0fWiAg3HeYgsw
O4QbP6+BqMr0aL92dM3gEIbuwNZ/cMUwOz4qjID8v4dx6G7PLCGBBgmKxGA1qhF8COg5/KwFpaSF
l4j+dYBGs8nC5VGVWpok+lhH3hCVsF1eFSDgAImwcRRFbFEIYahLDcU8lFLVNn4hgM5wVNp2TV0s
kXCMImV900mVtb1HeWamRTcqrrGkYnbE1TYLTdkf05rs58TpwXQAnCae35S21HOlVH1HDTVE+jYt
rb+rH4bv3Brf6NE8cMk9e1v3ErtD5Lrc6Fwa7THo6iKPNpGF2Rm/kQliGC1ngg4CzSpbYIqNKGRE
L6+v4nvm5YNHOdgXgTo3TbuffzPF/yVtKt/gDY3L/c3mL9SzPP2UaLPQDZwPvNHGE1VI2H6X1p6m
3TiMw76wAdJOKOB5A92yw8eJguCXOJ+mO0ueGn2amdYOm3h4JwwXNV+K3mosVWhH5W4hQ+wXmIIM
3PHXHj3TL6M6BXsFIvFCjUtmPM9sGa1eHZ0DY3VOWNcBfNz0YP+ESUPbmzw8UjSBu3ppkO8CDctP
Qw3LbNUX6+VB6lNfUtq4D8/EfChN+498pHRD03kaqwg2YvX7X35zjy1gsJgWKirMijkdsZkU22xa
yPW8iNP0XnEZrmfFmxSqX6Hcn5IvO00iG1pU9yUGqTUe45d+LFGevXhyRL4cdfQ3fS8UIDuBC1xt
4eccOulhzagXmVH8cSz0k4Qv7dm8dG8U+1wgYpZXF3HK+sOAW2QOQOBUNOj3YodqJ5XoTx1z8tmJ
KSwSUr9732MfDFuM0GipedT5p7RJCTPZv7wg3Aje1kFIUC2GnM5QH+jZMx2jv2KQCJqwPcyPYPi9
YM8jagYcWJMELLt3ZVBX+SB5q8DT2rE1wIIcYSMB6aiWcTEdzd5cbGhNQqfsUmo9gOeIP/DlZ/9r
VumQrbjOQtyc35rSo5lr9EQhTodkgMEC/ya1alL93UU1Mzt5KYhEnh52wUgNhSoERiwJbB00xCt1
2UVFYybko4Sfvb88D4sudXIJHr2ROh5HuDbYzVHzYEvXk9OAlTE+chjm3YObgiUH7mzeiJN5bgz2
ohX3zGsZZqWUth4TLE5gsu7L292GAJmoAOskfGXSP9WPCPThpLs6dnKQWTzxpKD76WbAdTbjFsDb
SWxR46QbVn33uDZ29WY0Efk3m/obadXdO2YvhL6W8MeoNNiTpZezynTb9NPPiXK1Kx8mD9EBZXzB
dlIzsngOQElZlZZnSgJtrPE7NiKqNx+AGxD+AqOoQVH/UgksWlprZKWk0ACY9awPQ6YEcWUU7+IC
OTc+yIVZ3wjQrRGtrfJI4yWfHeonMlKT7F+j87tnNsuHp93mnCv+xlzQSCYAx5/3g4fxtzw/VJWr
vt7JheVi5hxQ9XER7GHAwgD/rLewlKInEE2Yj2jf4X7yEIRfU7AkJTK8oWQ70H//KNo9uUmGtn/a
Be17jIj5wBUyEpQjnMH+ZzXH8neGsa5ZiPQOAqk8qQMYOalGVTidRUbeuMHTPxyUlcBQrniF0jo/
IBoWCOd+W4Ji6OlzQor5bfeE7D0BcfCwQjc/n4i7XoTgsl3vQd5xVH8yFhS4sujCmm1zXO79Tr8G
o3mw6ZXiEW3e+5NWExJWLfHkiI8P3m++fOsSh3cWNW/TK6yLq2CS5v2TE0BM2GWTiqdRVhXkeQIp
HIsPn0mdLOU0QcsISA2loHCg8WpBtytA+FQbtk+0D1dwQPrL+gmiI0WTlAiPYMlUhh1Xfnrc37cH
gH2B19SBYvZxJZTJ5UrMn77w4gSBLBOWIwt1X3EbQIxu1PsMKUKeyx4+LWBESDrMANPERHmw09an
C3hbYfWu433iYcvNK0dEjgUAkXjREtfamhnzhDsCbOjQId5GDH/nZeZvAnndzL6T+TkEBqn/Hqem
7xO1AcxSS6UFMUkbDeLCUNm06rjC2ojFlLr0gPWlzQz4fwWIUt8jQwBJSFLW/XCKoqML6Lzvm82W
//NffWOs7ORaeYtzlk0x5PUHB0h5zYv704iJ3fWM3DbsQsZgubDQoA/LSMasapILTjEt0IqJT7GY
ovbGCmq7JU+nL0Gw3UwXuEbYWFXTj80ZRujUoBvn5u47kMDPIN9GFWdKqU7KtG28dX+D1oscmUBh
m5j35fUntMd/Gba/GrZDCIYNr9Le+QOzGRQvlEnCuglHpeUn2/v7mdmO+YCWStR80JlXPUMY6Qi0
1r7z3DPpz1nrjhDnWOhAMvB+EmEaR4lXBiQID/CR0f/pt1hZE4FnQUl0BosjqfjCXnPgSCQiDDcy
QXqVhpYxcRZA9sxkX6ACuFtJHXa+/UQ1qHnxU7UNZNPMjH1DEdvGFPCK58mrwnPEG3yR9dFsWMDg
apsopmtAl6x/+m1f2QAePWV+9gwdeWxEZdYoKyNwMeFrWuAjPjDtSs2HOm5f9q1M1/3uc90ZHUui
j8B9dYxEViiUrCk3ZoViHm/I6BU2a4PmeCQ50M56/yJtIejwzhJegcLDmsC4/kzvf8sMcOOq931B
RNJrteY9jQex+wH1bAPF/eGqxziRLVgP1QowQXG+EwCYTlDaqqOlRFpkw+7QCyItwJRlMRGFbEsb
yKIaWcHL2nC2lKWGmSBBZ6C9NaNPI645ojxLHh19FjDBKrD5r+DmOxIT3jwtmepRjB75Q5aNYeVg
QYDsN09bXLFtqXZl/xNe/92Ti4SOF0MXc9UN5CLXVri2kHTrVPojfbcQMWbUVL3TzCpJMshCpiGM
qEWu8DyuyxwwI+2fun0wJ6yGWLrAHOztqgoFMnXZn608+SY3ZhFdoQmUt+f8An86Yf0T7iDwTM9A
opZp/fqvf3jR6bOIiDMsuabt7x4gUUNSNW1vJsJSvniFh1cBEugkjtMcsideytSH5o0Cq0YuPvMr
LQi8qwYPsg5UgepZ8e1QD88thDrHC5g5TEnODDaEwGPdnyzDN4zTFkBI0GDekV5ohJ1CoX5xgG+I
VTbk/BZmRGfCWCxEt3/Ow8qWqMvel/nznpeWj0IjdrwYvXB7VBTpc+JlnlLERE4xrOGiNHZZKvFM
anZgaPwk6/eDDRwctrIJP87CsbCbu1lJrcs580DBIY1+YM6U5VnXP3QZ0iggk949iaxWC8J/+rN0
rvUYwAPR6Aq/Q4d9PLSNhr4zGVtVicOMoDohpS18CICDPtD46ez/q6fp6MEj+Rs6odVPidezEx87
bCVItAWCLCbpIaxvVEMlnTuUoVnvGrYR46ZaLry8XjUor/+LIGcRup16Frtkx6PHf3Vv+2eQL1dD
K007iky9/v2c9PHcqHLzQ0NhTqZq2LMD5NCLQp6s+XSDufeAH8Eim29noK6yHLxpkgUbuO6A3xNw
NOFUC66aAP0gdMnzu2Q8rpNIlsT6SNCsJRc9k4ypVXOnK022qopwEdplBHej9+HDck9nYs1h6FiT
dvh2Y+N9QprXf67nnUI+GtT5xdqkmwtiSpp32A3vu0W/B5rbi2w1jBQ54g0TNZW5l0nmd834FXkU
4y53k4M+eWqoXj06MAryd5snAo3dvBpKIs+KUB5VRjrM6ayx3YlvMHzSz3FxE5AL3L689jyJjNvx
C9g/AhCaLwFlZHEAzv0eSfRNvB0YYKZ3c2wMbwyh66Jae2mLOS44AqirbQkdFzCbmXwEerAENy1w
sAsR4l3jiopuGjj64eqwInmPn6jWpz5ttrijanTJEBbsBv2I1aZeVDl0InLpNBCJw7WVFrBtuOo7
F8cuY7b+xp43uPlXGQydgP2A6ywwrlp2I+x59ew7U0RTrO9Hs2E2AQhAFne6/zLIdguv9X16erdx
y70SMAHsf/WO1K7wdH8/YoflretzbTka4WET24zPgiNtZUnOmjgLiBAnMiTcIeuzw+apOQpjSEB/
0gBJRK6Ux9helAQkJUBl948KagS3+SSnHpPYJmHPkCqFX0rMfzfsOv33yfnDRSScJoDXuOEta02x
9lIRV/LgpvcrDe4tpo4GQ8yKJMYohPnUgV0zdivvPhwaenitfkKqRlP2x7zmNCOuKoUVuV50OCuu
vI1WeNkWXf6+gksMin97qftRlzi8LfBtUEBEYZ1ZZa/2pXiJrtyFDvYL/TfjNNaLl0TguMJZRnE4
oe78ok0djRvCXYsKowBK8TBGzayVzDJGuRMWjUWEUXV1UVWj4WZy4wdoU84C5+30Qf5ufv/9H7Vy
u7diDTAT53lOQlvtM1PWbr7SQ5ZFvmOhrvMXYGxA91WZYiLD3Zs3d0DNqbQfHJPEfLzkX0BZ2oMW
I91pGht94aufnO/xNUrewqyBOPxve1LWsbPAbPrf4MWqjgjpP3fI1SH1ps/h8SFNuJtKObMyX4rk
1kfTHjDL3KsDeuldP7zf3FITtsOH+DFwgaTy86o4wEL7MZpmdgpp8gbzP9VyjktL6Vc1fyrQlsRZ
fytjXQtoKgkGIGzR/4n5P4hsHJ06KI5UliUu4B964l90JLw/D77BoNk7kDIVyqv33j1kuqyKQ56x
c9APHb/fOrNNiqEc1pZprXNQVXD0fcDVdMMDVEVmS0dCIgDb80GE22vj8dRtL/XDu1lBftm2yDZ4
YqJ+Kz9MVH5cfY8LCDx7q5WyMZm8PB9qggP1YaB8LOR2es4hgefu0pWfZsski0Bky64JS9xH9TwW
gUG8g8dFmZ5x6RU75ZzIYMd+UcbrOv3e9IhUWDeqilob3d99pzmIksACNJoXy9m8oraNyhc4d9Zb
vvuunZgd76ayYTLZBfHVVYV1ibqrNGBsmHCcPrJQzo4YX5huphsz6DZFJx/ovm6rcCLDaNK0hmxw
WhEvuYMCvbZz2s4WhDMwNsU+OepbKwm6gJg6Lo+s/dFztrbI4V6qhPhq+OjGme1sFuUItGMpE+sg
UBoPf3DU+5jmqSF6uJAvKW9b7Dw8Syqfx4jnNaYvTx2OxsX97K2WEu9aPQuvLOWnJvZAsTck1xSb
vK4DoiprQqaUa+Aj/piGry63LFW6d8XpEJUEHmxfQVQ0WeEJXdFp2Zx7L2kx9tI/PrrHZdFV8iiE
aNJ4ovkAvDNxKLcJPEKdR4bkT/Ud/CeRAjGcrVX5q2Csff34be3c7Na4mitJbccrU+HGdWbLxtyg
LNfVuqcjq31U/wi+u20eZb9qnHYa27hrseER5rLTzO1r6bLLAOQqF0ksWuwOsFKszEMw7xIfrT1P
OAwOmsaHDPD6eC0OP54x2RLhnT807abOsllUc6NpWMq9zyxuTyB3c8c35Ap5tZcjC9Mcqjh8hb2/
9+qD82wDO5j2my72UeDzPQIskS/zKf/MShG4sQA+R36aFGS+/KR/k2lWtnEpUYbNF3JU5XHAhjUn
QHUYXFktrYMjGCtzLsTEhjPoAbGHdU0zH1owSLkUzyyj5WIDX5p9QT29QfMX4z2i3g0cqtDG1coJ
pR4XM7aX8EIn0GkkfafosZFOAB8VNIlXji9SLr1p01nl5iVE4tfvo19BE6G68jUfB0OwFl13fBMB
gMcPtoguCc4QlsuSWde9ZRiL09I0rWnJ3vgZYAo+DbxzGqE6fREOAnB1I4opudvvL1nlTb1V1KZP
SbDL8zgawCgWF5RgKjZPsgdSJVJ6aB7it2ably+h24uxMC0ft3pBRpAa1YEd9htyDEb+UvVBSmiy
oWmsnFgH/URNXbs3jjlEkY4H49wVNQMYRXyJOC0tgK7mfIwksPXfh7RlXgOPBGaCyFWXSRWq7eIO
o7GDejzDGX+uSym73YN0FHlxNEI1UknuO0NTISqNCGsUWEKNIY0pEFbPAVDHGHVyn3pw/hzHgHEj
pArlisnVYc2xNhqsx+5o5wWm07VJpG39nnZL4zehcGFZr50BDKTktc5fDMBlwITmbL2BGvcpbO98
blv4fE2LKXvwnJvwP00eOVkuOVrJMb6vgIJl+Cjk6Bg+22Yo6TVcvOtDtheyCl8A5GvTicsr1+3Q
3ucTCxOo9Efx5sFWXFsT39xyX/fjol8zo6npNw5G6FLI4/dhsYnZ/Aqee9jCEzlmjlKzLuIUTtYM
Hp+eQC2tdcZ66RhfNl8dQTtiGqC4iKH4sUQN0MacN34QRjEuzqC8A7UpKkJS1tHRRzmVs2Pg96K0
mQAvQ24feqNheOmT+JCcHesExHBjvObD/kBTQddvD6ZYql3zCQDr0AOmwnldNaZ+y/0VTL2hUX2P
bLqZxh/YCTs/SgV8tVyhtI85T8BG8H1XEjFKOjXQ2/s6I/6tayPpCglHvVoDeJibYMu2b+aV0pR1
nfpmuS9BoeBX90JsWie7ok/2c1/L7EWcSa7DPcoFTMOlEVKVHW1QV/VbjPfkRh92fizb4QIazOw0
tyByunkrEE8r+g2Uc0De7JEmFwM25tA1vZRVE7fJ8dKYqWRUtlRxVsf7lB5NklPbTupLLsaxmr6Y
DEVyR44uxLo66kyHwJZO3yCRz5YXObNyedrQeQJkY5eDeH2wqy+70H4jmToM0cf0qrCx+y8Sa95/
mLQ9YGr2rE9uZILyiiikmGN+koh0zytAYl7HT6RZLepMrjYOpxHoCd/HT8l9oe8zp954Vc58I6x2
hBEKwZDUxod9CAU0RqZfQhO3+RMGZ8Oo+AbdvjjdOwMqjLvBZrUd2KtCpXADPMRo9Kx1MfnBUYPj
H82YHCTBj3z0tNQoslvhecMIE1hDzEqZQmd0lZrJVE18Hs17BYCj77YTiR5IPJMlb/FFAUK6zG1C
xgskCb4uO+DlfaRMYk0R1ecsXwagGpIfH0apefqWA8AOF0mBrnqZnx3mdgAntUjTCqgwjws75iFI
tIKVCkt+J0bl/FH86oK9FaAW9NIopc4bmQk8uG8SKHPtuzNjXl78SJCMhsWJgd2M1NHei8YJgY7e
rZJiBOZhLwpMR+N7BDjuY4kLLDug0ivyKH6f9voXxjgGUulId7oCOz9ofUdVOERHbuMDrhJhkiGQ
6VYav8nxMlZsuZbIpkQy3IJnpP3NXDl2zAQaRKPYuykUVW4XVWH+YAINTyxEaZiw8n4H9fYqvWZq
MR4fpJW/CBSU79Q5Pbt7dmwKovCMsAoU/PcZrqxIj3eFvb0zf/w83otdn+D4UNXIfKk5XvQfuc20
7PSfHQT6Bj7CIr+VA5bmtcrmxRlhpdjHyXjWrpmV0f/IwkG/q05rWRtaXBOmvEdC5KvoL6MUU5hB
Er3B2wwstTI5hvSCTAbkih+YAAWatckJ+uyB/UhcVbTQ6EnYJT/F4gUrkrl1vamV29F9NSpsUvW/
eJYeUG4X4ewITVQ7ZgSFQWpRB4F4m/DgAR09N0I30VFNbFkKviZiCp+4q1BFvVJN+9CZcGHaY8so
qx7fHXrFluUEJIhZ5dPPcUwA4FArNx6TWSmxsrh0JA3W/bl5ubxt1/OcarL4dEMSxfPsCqYyMRZP
L09oIpPovm51GLlTuiv01SbmgNr8iDSxa0ukSBpi9oKso6GW8MQUOTBeSts+HChubGCPe+f/HX+L
WF0IgyM+rRxI1lqmjMFbOrkt0DrBkW+QXvKxJ8+NexzqXYzIdihfNup6EkWMeHhlepDurs3lD+VQ
1nEfCyMBut/7kDn2OTTSm0/RCEqd7rPD0FszPk+CdriVHUqiDCmMnLB7OOEvPlBTDL7JRTdsjzff
tsrL8xChzxMusuB0NwNccfc3rklAFaZh3jGuAm8BMeZbp5JGfQUFaZMwoP7XXwh2fbfsSYpoDWE0
q3Gf5G96e0Y4QnqykcRIH+G91ThRG6LWSK4lqVIiJZ0LY7ZPVqydjkOb1jYP+mDbDiLzx8lxMnEB
sUkC/YgSgV0QoGZkBgVlHds21pV88hAJWKqFDMN/p4z9L3eQnnumwz5xBgwVRhG0xhhIBV+JY2iY
zl6OW6XWYK2isiK3Aa/fAMHSYazxN+U33vniFGBzMC5zd75OKFhEKd6zPsBTMXYdCMRqLlH6RA93
/IEAYpnVXC+6auoIRE6qejPlNYNChHZjOXoc6+uAqSzgZrCgBCUJ7DFQ6Ch5xlGFi8b2Sqg3J7nT
TubGUrq9fFypB9xNvMh1Ju/tQoH6eLAvxUE1+KrGa73p5GZBAy66gjfcC5IboZ0KBiYVFSk04xlH
MdIOYMMhTVI/7NnsZcStEyQ8HILlaz2zzAb0fbrB+fga5iLFZBh02Wj5CatDH60mI/FTJv89Ikg1
DRGHq6e/M0LeuoklRB/g+ePI3ELpP/RXHCWHVf6OjJv/jGXM+E1Jb66HTlSi7yZD9o8ljTiXg/Gm
2IoiX+8tY+/uCu5LoxNR8FnRZEuGEl/eo0RGALoFKjpncqCcxZ1M7m1WkPTahuT0ddlzi9ZBUo8u
VxwLr6hGZ/XTOByjVXuWcgfYHQV30a+sdAX8WMBCYyz96cHOkZXBvQAHfTpj5Qpduy0U0asa8FHI
MEM+6MBsFB6wVmBl6J4dZYQlPL/PLrlODn8BJCqhYLPaTHiXCMe39ynO4OklmQRphDEtpdseTHt4
qf/YMo9jEfqJTIxs0JM+zA5ht/NnW1zPeNB9CiMhpPYJgXJO/z/WWhobKJ8ao3nsDxRQxIpqZEIq
VQjE5VFYuzbd4buwjDDz0Vgf7s5ionwsK5Js0UQfGGdym0KPauHHV+I2wr96YNELVX30Mf6GGCee
R6pCoMx6dNDrupUqrqrlsCTgqTffX81dwNjES2zMxc//rRpDVLdvV9n2RkQjbCY3sdOp4a/2f06C
vXcVejT0oXaDbCL5RDHOTT43OlMY6Z0exFTSqokQB0IcvXKFGEp3vZY8LwgFgo3WRjO8fK1ov7J2
9aOrEqgRQ8KSl4x+SELRA9GtthkDQFnotJn0vEF3cLFGzb9mTUKljtpj/WU/uEWNebtwGHAUp0Jc
6loTJovGEai/4DpQ6oIzoGGz/rnM0/pCgWuqR7BKkMgHB9qwbzmR7cwcD8dzxA1anYTzu5kZ5F1y
wB59GqkMtd9QGwzjNBwRIVDrgoBDTygp32uOORgfPAQteQEZM9T5/nHLNSQW9G2UxDtYxO/yXxzA
Gn8Wgm3dpzTJdChvQEQjV/3XbUXJDgnki/r1/sw7JEG8RXEbe/EyWSYoM1Xw+pcKeeb4xyq57sqa
uszXo8BmWWnT0KhqKBRBX+yYak5kjjhb/8S3m9YCTNaAW2gZ80ryZttwhP61BFIRAdIFN//vKgu6
BnIWgKxy1pBy9oIQmra+maqgKCFaGI0Zl7iFgwg096ESc1YLUX4NbMb63pzFytlqq/omq8XsToDf
exHM3srKzGXwMbeEQUfgbRndoj4rAi2bajeKEEEC9tbPQFJWReCPucufVB9/489eJfTQioZmTkVj
RQ7ZNAP9Xat3ML/GbfBtUQbfXzRAaFMZlCGarTKB2XsDSd0B9LGAFHcZ7pKG4eiGLzG2Q2fymPA3
zZwJ+dbC4P2DvUIhkyy1SkstNkpYRZE4+rmp7FGXfCI7e8qfwoaEQRPO3DzQSqlkzZrzIQhP1lb5
BpaXCUqUSFqZw4nogrixUVPz8CrZZDk2A1QA/BeYj9lUDnrPjy+02K2iXaZI5c71lW3IstUky4Yx
OWQlKBXcZtCZzQdZL3dbYqmoSAD72PB9GpvM0nZyYvmo9Sfbi4o0NmkDmuURSNg7lE3MakcDjq0F
JhwPxImwJVI/JV2Qi9AKJhJcPkEfYdunslgtCWMIc1M+jm/OvaJGJNOqNVbC3Vt18k5MhNydIPd0
tXyV1/GFPTri3Ep1h5vpYdlfUkVIT0IvIRluhl1TgkW5y2vu9YH0z8TTEQLqdy1TP+hImKYTmz8A
Bzqpbo93IgPsU6ZyOTPvz6Bxb7I1OfYwe+8U5RrVNaQblBWFH4H/Nd6q8/4KUArGfYIMhc5kdua+
r4gLefsszHSkKrbQ0t16UISoIZ185dt0DAoc0FmC3ZwgkuFj0uIG+pCcWzb2DGAa+xPnU6xlRS1T
v070LvpZo9C39G/O7YFKnP0MJhn7PR8H3HCnu8SuoF0ac+AJ2t+E30Hwb1g1P07SvU2h6ZedeGGL
+jvD/QU0irfFQ6PEj8Gs3Q7vApESKFDDsL+ZzWeiNwLApGQJ4BlNQIKpC5Todst+/Fa15Y4tWjvZ
TXroZE3V43z5h4BGj2YJaHz5L9RP0kvZripoMRLCWl4S+hSLI2ZFcTrzVP8VG/3ZEu1IsnNaHYLH
JQjhzJQ9cHkyfb6BCrxSgulxAo9KELsKrEF37DXWZOzm6qPDqQ2nKs3nDrl/uVQX1ViNRVcESi2O
PfXCvGilAIggbSUQSW0ymQiFyjlEDyNhgfACEZtmD1uzNZPzX0LU/G/iWPpiMn+oQ43y3QP0fpt0
lSr8rWVhyzsCHgK5JERPklST15rGOLJJUXWaY3FYjm4OqFdGmFBNp+RzuQkSmSBDObgTDMstBxum
EKINu4fMJw2q9lvtiQLO+jGkldEVxIxfY1r4e3XMpkdL7SDgLta8rBRaJOrHM5yYlXH8Ekf0aZHX
HYCEneoab6A2nt7eLtdzvkfAwtxUH70ZjUT2KrZezcnhFv1VogC+4RijO0KkAleR2UwARJgYxKNX
HK3jOJD9pXpN63l91MGo0wwAKJNY8IQlRFTeZizGBxSwjb1Wv3+mLG2bDKd/UVcCnWeJvybrWRER
l7mwS/cC0z2TCJXk9N5dmQn4sBM5vP0zjiSh/I6bPYW2NKPEXVTHhDREilwoz2V/szzwORl7Yoyz
40V55RccVapCGohLyoURIDdNEZiyZCO2xcglHeWJv1ocuJCzWyq3ZPencwxwTYKxmXDonI+m320s
XhJsJpIy+N9AlP5rhdKBRbaXVcmnFSqTYpNd1sNpdr93Zp+zTB5W3gnntbwMD0dFs9uaBVAeF6hA
UIH5LhWfoe4yJSBDc8HnAVzsYZuWgbbP0vwNmXg+68VjnoBpWHnu8WkOoXo8m+N2fBazvsqPI0mw
jmvYr9IhAvQjhGa/YyL+lwHD3SkAze4Q9H9uyEGHAwZNjGh1mpsfR6VUzOX0lz1qKSf2brZX+90/
4Arugf7B6GwtadRkdLer9pAjsAoV3ySjx7R7xd1ZojebipN0klTSM5bIyRcX8cwMoRrGAakXnu6S
hrYtnW+FhbRCkxh+T8a/yLW198/vobXqlTcSvSZ+ckqXSnqy/8NMt0eAGi3p3AnzH+n9k+PjLkpg
q6RFcRmg67DgzKs6qSA+/4iM8gPgO6LYkbqkCVq75RntQK/nmZNNi3qslyZ8AmVeMFw+1xWLTZgU
Sbq0ZVZqN6OK1Cy4W1pPGRIqum0FEhG+CKJFpo2uWE5e3CMUTi35ZRAexjEbXohiDEjlsxQoQqrG
d8hyYJvzWdEBLm1iqACQzVwBVwVHvJyTN5xUqrKFSIzge7QXL57QLKlHkneqhopeqoKF+DjMcW0M
y08EsmXSLIpoLLndRxQi4WovAeDh4zkAoGlkCFBPOCMY1/hEIDiZQFcH/69561FgUNhHuVWFXSDO
72e1iSVSDwpud/x4ajvfM7ee4HMzw7liVmG3SPt1OvwUK06comROEI5ezM9WTCy9uBSyDKcjAmM9
uhOvxyT8QkmoWYMP0n2/etiP1I0hHVxNwUOFWoAfEYGGNSAPKXIL4Ew+F6S7Zzk4v0bDR7S/dF05
oj8GbX7j4hxijyxKWGSs0NIpvSClnuRgufmafSSC4Rkhcq3/cHbl+5UqcbHqDP7+YvMmojDTau9j
EfztT2T8jtstcpHCH3K2ZomoZL1qzkBIQmwNb/FxcnXqzuYa8Spdxk8WplYW8FZx+4mfRL4YlLaZ
Lw/ma4Chvuuqq1NjiE15A/OsW5x37Sdv0DO0c49o554QvwEl4KQCpCKJ+vDrGiwd3Mod6R1YdZXx
R99i6riDFA6XwQYYNuio6qvAdJI1AMaZ8oNKudcT6h5SWifve4jwQxDakDSWXdhvY5LLY1h6lo8g
Bvtr/ZKeiUhPdX/jyRWOEEc8YFfLDJ7O7T9bB+X2VH1mXsY9Wp6ZKSimWLrOZ+53kxnJNZny329x
iNVaRcA8Hq5+rviOm1J3z/j3vngVvAi7DOcuIvcJEP3hrToyg6p57XEB32glI+1gSsMtN6Uc72O+
c4xlM+DWbFYpIsiz5ZOcbs/uXJPonm6vmNbSu1jAJi0+ziqhbK5BErSl36Rz165kdt51MI5lLWDJ
83pzfwiQvDQdYpvX3pFMKL6ZDjWAdBE0uZnPUP75bdZ7kz79EcPFk+OOjLoETU1/JesdnWMxgLqQ
FlyBr88WiPDaQOWApFRWwoha3IuJ9CrSHxRUCIvnVNA2dqrugOynpIbok8Gs7s1imgrDX/5vXrOh
+jhbY197mU/EekabxSoI+iz1ACdBJ7AuyvkKwJ3Ujv05C3AZthcFey8IqAl+CQhf4td0DHoM2dbS
LSSPsSN2HAhWpcoIs8bdHeLj69h1ZAw74i7gMO2KJ6aykXfNdRcjg3sblZZ4Z60rQNE8dlOP5YNr
AxmaC8vhmWD1K9IA7FT9uCxPX0B3EiDpkDL3S5oVt+gl1uPDltRkjBZgMDoTqEd8E6MvFBBnsgkj
A/nYgIeFinrFy9HAQQOGXTM3ircV5u7IG8TvWJ9y9u91fbl0nlEOhiD/rpjquJKScV9vMpb0kBuc
BWpPdyUbe0WCcxGVbUVpWFB/qI1zbqMbsEtv1RAKTj4PSVdUyNOaCIxx3VPDBtBxj8u2Bn7yTZbg
ghyiiPeKvmnQqTLoKqUCEnDmcRYQFAaAa9zOTGKHlHogwQmruf+Gigay8I31em80+HrNrQgqw9nY
ufEtUN9cHrD3S8tzoEgrmlY7oxFSxChKrrmFW8H2d3tasuYlYWuTSBw1WZoMspiVfRq455IlWhgk
CBeXYLjDFmzCtESN7+ZkqJuU4WyvoYBMYx1j+Dark7TqrpYvKARdykJvuD/ZxoMTM6OskpVeTZUU
gNqkgQjOpsr+PaWfCrKflRx1EpqDlIYAzWL3JoOzEce1yu45StxAOkdWSvM22+fw6oY8jdVc1S8i
sQNJRH85ySutLyIBPjW17eeyrSYaTTJ68of2QuMark/trEel8v+mO4OqQLCcyR73EKElFhMhbUlw
jrSifUOQN6AxrG6FUBonVFp2dhWpWyC6fQdB096+3jf6gRr9BhkkMmFwnjN9tbMQWtWFEWzCIdMe
mBFAdKJ4nGcYh2piWW+3wLzREHvVtCFk3jC/uBqMWzIWvofCs0Q3Cip4rg894oWWHH/oNvjcFAmc
SiqlSJ4WSk3NbkR7VpEVaqVJwP363Pwh1wG6eKgbfAoQEVEGv3yZyBA6v7R+kw/H2NwEHZ/i3eKJ
1dJ57Bs/GAfFO6GA0Gy3aICQQ96aBypWyOG7em+fu3umrwP+3LsH42AH7dNx3BZzJDv66bEJqgr9
fsSF2JM/RtAjMap5Q+UeEkSqYyJFff6HLhJ1UKAa8CVarWgG39MGaAvy88UI+22g7o/XJMyb/9DO
+N4bYE4UDI46nMRNHNRhqeDJJw50u7usHHc9vrbfrY0/gJKw9I0moShxYTUtW/ZukzPgKf00XoWP
cMoQRYBSW2/7eeaNNT6dbHQ81WkcO7uiKfNVXAyUMQHZkori6FZM0gMcN0HMPVUn9IHI2raCbltm
pVlIsSrBatY+xCCiYwV3UZW0b4D/jy8DLSsN+rKmDXxEC2huu3zC1buHMgaie8NOH5E9QDKlQUWM
GW5FMjahdI7Bj0jSEC+ca/uDYmn7MG5qmeT4W5GwKiaa9Kv2v3Hqqx2NIZ3yW+hpjTrVbRyfxdHf
tdx6fGpNYtV0oagYtFGF9LZnojCneF3tdFUOO4eF+jiqsWPXmZ63zQ5RdIMN3riLVNrTkyOmYGtA
3AVR5PdZrmSqIv+yARVpjcqg8jouqWpepOw9tBsTLapVHTCPEoXZqIj3lUgfnTZwEoJKzG8s+oOZ
BwRmabQY0ObJm49OJIJJkUaxTALMI+LJ34JgJdf27aGsXZtWs+60U/Ub2nGFKvlLFNmI3l8dScdi
iP/he2L+rDMXIXEgyzHoBiJH7njKH11XZykwUWvAbe3Vjlxmr5eMMT1AN6zb9Z3SiMf5uU5UbhFD
QzA83FvmOw9oUK1lU4A8QFymi8qZc60XYEaoHs34KECjUUZh+tIsVO5bKmXxbpSOvGr/kMUJ420D
m1Vv90FtwPfS/jyqJyndK0ifGWVfAK2H8BioR6RsRDJOjQdatUNm2dN7sU2dhSQEOfw3+GwgMiE4
tBW+qJfYzTOD/mJ24aq4zrBm3Y2+szngBL2CXEVlDB9tZGF97FeFv9VhLWDNupfJ91O9EgZ+ADsf
oJpAt4lHsyIAkT02Pbsl5DQztWBMSUzIb2uTzqNiUzZ5LE3Ka5ED2qHwqTpieSQz/UQAMI/YL5rK
4TkfS/DWAAkokLqMEErHElM1RIh7CUAyp3QWU+TWtQIRoNo1fvBFctGW9Acwo4uBw762VjaHRzId
CZ+Q1PE0E7sWfgQABzws33Pe0LBwMZ7K8rTUEg5VKeAMjs9PhGq1MjnGAABgzPgGcg9G7tRqRgG5
LLWmLoOX+TG3UKHm/SNamb9ruBTAVvhZ7+GK7k6f2TIazIE5Ilk5FJNbDn9msxo1fJDljqt9zO+k
Exfl9N/bCmNx0n/p7ogNtBt1TRtpfvOwA8JY+ljnq3+BZ6BzS93wLtpHUsWdmkkuFIeOYm4YQ+dG
MUFlMUUyt/jNG9XEc6vfo+89N0wwUvAnBQiqebCQKQn1iUrstNPfPdNJsoU8b7kruU65ZlyktK1O
Lp7hfMSjIXPkKBwyklO//4RSTz4qkBBLsU5VJ4NmBangym84fzPvz8kZ3b/l9xy+9DbbNjD+d3ql
j+hrTf9FisNsg96fHQ/wqornys0S/LKULripEsUyrUG/5aVdBsU8wbpMSMonc2P0vV/5y7A1TSbD
Esh6hXYXSeU/haXRu3wl3ljnN0T29sTNLbnBDEuAjwvuMrXFh5FH0CYj3Z4i5EkHZbp0+12Nj/tr
/roBTLHrmvzQaD5vf0MfLdzu2GCe7UU/6y3jP/jZ7VpyOQBovwlg2OQlpPnPUM2p6wNPmfSsudm2
K400xPfoXq6/hPHP3WFd7N4cNygrT+14f5nPxd7ldajgWfhvrwv2P/5OR6Dk53+Wks55Zayd/s79
jwj1v85ubVmvwJkgS0s3vjGehdlpJH37C75EJl1o0583m+OK8+W1AeHVoaB2NrCCfDs8gdjDFcUX
mshR4vAGHjr7QmG787qRuTKW6ugbd6uu3KO//p0Pe18NmfZTZQUv4AX3Y4kMYQ7Qml/E8JL2btSd
OCCupK6JafFlQ9Xr/0CEZlrC6qUaTW6lfCVqbjGyEyqbClH1c0D8xncDY9hIug9YexZWmPnZziOx
1afzGu+KtXFdaqKbQqX1VdOFQ7vRR8eWNU6PKt7q3Dx5v6IR7feSlAgFubbHVGevI4CJwQWiDugk
tiyAXiCKDIO6QpOarpnWqk8CZ2GNqec/JkEXay3SCtm36koMkSQe7TEKbClktQwfpYAjfr3vr077
dKV6h8+4AzXYJnIK7V1dxjtNcEPyey+dRzdE2h8k/5ZvghQn4P1IVLQvdl9MRAwHweP/i+wFUPto
2cdXS0xS7EZrFuHg9nfyJLMAb/O1SI/s0b7UClKuD82axtCCWkOFE/1FzmUomLYyzOD+bsm3Xg3C
BbgXO6tETHlxVASD6Z+HKQDnnzEhQWXSr502wBFNvQW6BfxQjCcz2jkwsvByuxMeA0/ttfBOTZlF
hxnbAS8yWVYY5KA76N2s+0RHRzWZBOpY4GgPPEYVkavPXU5HnQ8u9LA+mDb7SzsvDUGM9sdOdDyN
orjXeWWz8DOgozZlePMOUcr3l7llIHqkP5T9bvwPj0ItdtDsO9RgoWR0XXohGO3yvuwcuOQPfCSR
AKOSdAIZM6gn4vAATNzHgQtU/N+VCj+Bl33zgdWizmCfrOUEsQbylv8nifkubhxE9x3XBVz9ds+Q
D3yE7JfG7ExU1QwBtobIchK6vgxXDCVluLy9dTQRtkrWHwPfMKkmJm+wzMHXD5iGVNEFqxWSx8pO
J3abWhjLr10W+r9QAmhZjbUCAnE4CjsHvut9voC3k30JkFisEVNfGhYCSL8KL6DnT+XY/SCOxJ6e
8RhHaMT4qXIglFtL/pJs3dKleE87OETVxGe6pXOGkFNRw0FcYqm9D35IYS/y1JZuvhdHAsFH9PBg
6kiKMk6TZwn5U1VXmq0Giz83z+7FXbHw+Ar5MvF0tqk7uJSf8MgsXsH9Yc0sryzMcyBakrurERCs
W7IZbU74X6JsdpYnY/ZxAA6MWOEDsJDk0m8kWxGwJm4Eeu2P4tBc6OS/RTwP8YecXcJmq2r+kRK6
NMP7Rg8cikW70XITeUkzdshUuy+bO79OaVNCiSIO/Y2zioWHvDN0AyhLkKQdU9cANr7bIJvykEpZ
p5bZWJZd+P4U3iJPnzkfbx4xcNiFKDw9C9Khvtii6g9olY/PSH+1qUI65k4AmxbvOmbPkbHIBcYr
24nINtdXsgf5vxTgtimrCau1Fi9qFbiQV5fHSSrBC1hYGAKpdHYRwCgYAwykGvCmfrldOHIxM9CN
5s2U25Qkxi+v4qd3GFkjnhGlVDA5E7fSP73GK/+J5KY90OCdBdqOqSFl38qDgkffs95bpG0bnfLz
5ER1k/DbF5Q/a8lcuXBbyUYZ/96hm3Dhyva4/BPaN/F0gF5nS/rHQRSwNza8Ea4/VfcjpuK6SQaU
AiUQaVpVPT7WL08V7ruCBG7kbHHkXEizwWn2824eAOio7x0gvG3PcbVGR54HiddGbOvxr9kxgOWS
+it/cN0HS09EWBgrF0DXwOhINS0eR8ri58QtE+oSefpUtVwIm/pOXsbAoAWjk2F9HlauIby2phBg
hdbaJJigYzS4T5KHt08NBHzep6oXWXrmzwb9Vy1RdnpMs0bKXCw+ZxZjsOS01rLa4xtz6C1k5mjr
UIcNKIpX6sXNWaKvnUTNAjsUtiWgqS6Z2PXgBmNsQhAxfIk+qAMqbgyOB7XEQxC7VVl18QwkZFf6
zNkf0PSqs6kQ4a6idB0sYCI7/YNTRxtB/fsW6Rhs5m5iRrsvlXEBtHvns4cW0t4CHbtoB/PXIfMM
ZTk7grY4WtWfhFBNMDOBE6DR2yz1s+bqBcR6I9K08apfSF+i1jbNO0RdMqisCLVbSGmMLiNjXs1p
Zr51Sw4GdT5QTtLHpDtCzxxHfbMWT27dypSdVgSVbZR1dQ5GC1qq1MoWdGGrbxL++cnlhdZcqnnX
k/b9ridtf+wcc+OQEDK000SUqkNxjMOnm7txzHEBVhZ4+0A3kZBJFr9hJzpaOVfuvvPbZrCK33+R
ZthkFzEM0Q9jvjBgfUXxxngfjtwvc5/k9unUTOCv4gbsYmsVStub+Nmx2xQoUUszV+FAQarEm361
oDi938S1bNnlyuqJIII2RlNbKigKkLUGNRyY2pdvQMqOCF8eMaS1cbPRagFZn2AMwVQSO/ccUd8M
1Pqe5vIN2795CZMKgT1cek4q3M4+o7glemD1IGXcEfNLJyK3jtLaCYYN90u6oBIQFc5Wp1IVpznV
AbxbsirESG6FK7nrmDtH5eKnJl6Y1bscfuHXW5htb93ZrWcJsaI5YnqVNaUvu5HioiPY+LR147+S
ZKy8RZJyRI5RDny9nmbzEPOjokPYQpSaESQebJLWb7sKhIrB1naqzUUhLHvVvmBaStDq2mEs6ql8
YEewa2W1zQF8VYduChpfVpMEVV0dqBRTKewyvBsjO4/H5TQ1zlh1jxuUC4qe91z0BY3YJs03u1Nt
kD+6H98vxYCNpFedsa3bMQMjlaMXz3KqYqTV8mGmZpbJFTJZWmEgoFMaDWr/XWFvDpuMlVrnNhQZ
SIL+jIzq+rJNiqNJ/oV81KAf/mFymNbvGcWq9T7GZXOLcAg2AbqtaE7aVmv6IPisUd93jQGJ2hYh
nJpDVNhGDCxPXOhONqvneI3TsnfivL80K+uRuwr71FTGdEq8QJzffqEy8MVNqlS8BYi2juLc+HhD
VxfpUQbx9O9VBpFx3iLePPT8rOOkt/2WsrQ/6+ley/lG6jj3BxTSPi1G/h63LXiKrxOd/q6j0RpA
XFzTi9XlAGn9cb21cuVcJancOchPgO1iPRq/OvYcXZyQdEqqK9E7/iEtZQcakCHv6nWEmZ5YoZm4
a5iUV87/R4D/4D5/nLvRwWaCs7Sj6kQjOCK+mn3lljK+EBih8lAWqra2VTbKlWS23tBw3v4mtt7Q
Zq5fos+Qmfv8hdFaQtzro1j6Bmx0LCe9U6wz9gtLrPZckHKS+37gH/qdC3WryNJ0EPKOOeP7sJEM
e9EzVc4kbkE2nQnRKnIWZ4LZpLczTjdz8/BnM8ZdUHf8Jhm8ruCLeZNyQIdPCABAUF5BVD3Ddnv5
JWReQY4Cvh/b4RZzTiaylH6XdXeEWBcBEA8siAdGyb8LxWku34quNRqaPjV/rJOTp4krO7qzmbZi
j0j5YpZcnf48k+TCpNTDYDgINp6vIJOF+IQmxk2CVn4NOkA5S537wuSpyqBssr6FsJBzeVOmuXho
4Yc+VLLsn1lhlzf5jkHl0cpZdZ9jjWCUD6vW1H54ZlHIacXMrjgS6aLx2C5p3e5g+VxmT4JHG80l
36nWxbnQ254RyR/HeJF1W2kc+vB4jPagjSHEveg20LISeJkkdckRKKym1Q22OR+b9hoV645B3J6Y
DtZFqheX0v/xr533u4e/R4dcGCB3ikQKSQhb7kKNQbvz/zoyNx5b1LijTeA9rCRptvYyk2xwMoJJ
WDOyMRruh/cvfafnnSxMwgOHDqL5IyTkgSe07qfv+CiBwxRcbE1Xpbe9PbHxVuSqTJ/iZwEpyuAm
7fPNXmXIWHmfmWJP9IOuUWxwin0cRUX2slD1FSTgSWuA7h3ogLWVEWuUOkotRHzaZcNiezJ9AMLl
F/h6WTeISnq5LZBVWwmGBsvRRnWLEukO12Gtbm57XkRcxJYdrCcykUPFtMvgCf9yAupR0SuwbGXE
K4242oxl47y+m+ry3Tv4DiN1WIZwI4rPS0VNM98tNQT5ZaHn23xJBohcL+Q0eRXDbo9aZOFkCPkB
MLUUsrABC6iqCebBgwdsl7NlHbJ4rRns14XdNLNyG3AvitejW+b3BGPbQ6FuCfzV1PzxJfL2+Jyb
8QgL0jCjYOdTR+dQIP77MRajCRzhNRU0snMl/CIRpj+o+TG0H3KkL4vC0YbeWcS0g+AaAmAfVloP
NPeEYojs/eWwWmpqHN/WFxEHAbSWVPyf64nErBeTlHZI+/vcdQS0SUD9YNPQ84zZaARVginU9WtM
O49E4gZytb4PXOARWLdEzpUZf0/2RKkNwLiTPRiGHRFsOI677IYZQj5ojKz7MSxkS/WcDSYu8Zr9
yJPQEqPS9jYgRBL6uiq1+NV6PhEC5afTC2SBOlfgo1//4/gma/EKFNjp6zQWzLRCHNFOncKK7+Eb
MZGmBQ4UAuc+rSI4Rbyj4ncUWYxxWtFJtssIXftivPSRraUgQKZh/zrZFpe5170oqbN5eBPKyRXk
35wtH7V67l1PXi4ruGgmjusX/qfB2uX95nqChk/hCMk1klK/gyblNUyp/azRBQzaEXG2LbPH/D17
MgSR5AuGoXxCUwUOW9P4Dzd33Zqjcx2/E0QANq7Xrj5RTgHQ0mBKDoznsu5TzJCt+RUlIUM9Zcz9
sW4aBhgyN2DX4o5egce9aAWCc+kdR/tfQOhmrPNawAxooGoNS3QVSiLc0GNZZP6xniXK/Hfo6iPG
m8zQ8f62EzBVPRBWcxuFsbIE2166UXFp/RbkxLj6JI1Im12Y8FVBaMngxPseFkJHRihqIv3WHhlH
urZDZNzhHImjBIi18f6Wt+1VpC9DBfgqRRGsNAmE++RJ52HvpTOELPRHRf3VGg6G3ZfXfpbywvdG
gCS/J4UhH+r1db8+sNL9g5/iyooVIYzXbrSvOJLkRv5RBY0PNC4EviE9gLWTaWkEDOrbcEv4uH3M
0uRQcrH6RqEhy4T2omYbxf5f2iXgPvkGAtTQzBjVlqXwwB3p4XxG3QNLP1I1dv3gznapU+vew5Ut
pMx249qK+plprEFuldlJv3H8MnS72HN19W621ukf42eqlZKfctwS2a2qtinl1mD7QodVmxfTm1Xz
u1073EeaUOVcDYXbI+sudUrqtOwQEht43utIQ7XUQ2Ogah7qyWaCMwqxvYEPBKCrZ6QB3+dWqK/n
g8ksR2G/scEcQ3dTd75NXdbYxuupM9FsQ/lN8C29VqCi+TLsjrbloHTSfNXz3047Y2dLan75aTU9
z2xlE0yzToC6emWKwT5SYjQIoc3WzpMEUHKWi2nKKuZx5AleOuKKxMWej0/MAfPL6x9fi6SoCIHt
0nfiTYHwu9XEIolvKwAOT8jCzKeO6zk6GVSLVz4Vm6c4mQihrwh9lD69ncWfqWxmORJvtd79mlGc
APDuivPIzdc1EQw50sDXpFV05K4A0Ksj+RX0D3LNXv+TQgvQaT2QwfCNnSht1Wx9eGSgqgfMdNXH
m8CaoTDkLQYBQGmiHaXJQ4Z0E2ZBRifvUMVyX33zswj0oN+3yOX9C9OlRUMZR1Z6+cdC/aEUQQJ0
WwLs4OyuaEoEATSKDZrg8BLU2UBXY7ha0TeqCc0ZjjHtgDbJkS3dLxjoFsrQoyNjtHjntq/0flNU
+gtpBQkir+bEKBW0e4UxjPRAb7tN0YJVf0SWCEmaNDk1Xwsp4qAvdseji27EidbePzqZ+TRU5pD8
zC6ul7xcu11pBmbZu+yAvhL6RkMZgkYksiQEG0cVa+5dxFWHxjspXn3HnDXLM8kR3SK5n0auSeIv
wKLid3duNhgiO9hKzjDNkhgBs71PXyecN6Ad7hG5vRTcTLh4neBMxtRwifX6NywBii1Wzl0H91JU
mVuQJkyGdzql0wflISe+fDIKBu22KQBiSMIbMRGIAtLwYZPSD54OnFdg/dvP1VY4bEp3lJq7QU46
xARKvUbT47HxQOsfGU3akM1H4s2GBlnP0PlQmX+TTiXKMu1vgBtZy5SDwlUC8pURDyfCyigJFsjk
4NxYqQvjn0O+/n9T/1oL8lNiKRTrjfO/ubKUQLtaT4kFEvI34vGbzJTPPRchOat86Me0xLrcxSfF
ExIKO34z1uLukBTNkRQM4jwbI/1zEgR6mGCG5kawBhQeJEqdF2utlcXqEo68DkswXr9T+YZbqccT
bs4zDQUlLNgWMDn9UVz3fHXiY0h88vQeYBoF+VjZrmnBX6CgjxsZihBtMqQfHvkIrEIRb+9nviY2
tjPf0H+wwlalZYPbfwjKdGjostKyg5rJe9yEsFXzL+7F3hRMZPQuX0Ybe5bLG5we5iTAHKUf+g7n
rRAVbWjIWgUl4iq8yd5r+PIchinL8xT9G16/tDiSRL9kPPDnkulGnKlKFAbZxIspVfRL9Hy0GZIF
/P+aPLvnPIIE16tCQQDC5dM5oqxeXxkCpY/P0sZuR7S7yjsGRMVNAJFOtzHdPeDyQWoTKcf2Lqpp
wcrM+O5cNHUfIXBSD+gNEODYQV+0Ysk3G2jaxMtbvuQSmdbj6CoafnVtTG4OYe4zstU4xaX8EIJy
flKtj+r2h/p92RR5exNtnyXBAGSZWcOkOdBmC4tdlNFFviiTqlpZR3TO5soJKhLA66wJPmGSyZKn
85+w2rGFxwXA0Pgq7M9kZn3Hv5yBsFeOMLZKhOwu+fSF/6NExnS72JNrQEsoeD5I4flX2bxpfyFK
Tt6JKqB2W5Dk7SrjwtDGtQpyjIm8ui3cbEaRV0CXFFoIq7l3QxM9Fy5uXHYDfG1YUCZiI8L1WjuC
TIybe3BiFhCUvhF7/ivnS/XXRz0Ah0UnCdaSYpXXrTRwD+VrU4z8ho+OmX4CGC4oIT5ZKPT7Eitq
2SnNdToBrNs/7w2G4n5nfX8swxOkUIDgPMVbnxb2KtYxWper9HqP0oB8xO8DWVFt4S4XWkzjMTOk
S1jmcx1G0l1SGHMt4+y1kJqMn2Uvad3t28R68rBuNkosxxoFpjDXxWJ4mERUQniZ6FkazbCpbqN/
4SP68hpIn0z10/PuOGv75mqpylr5EnTtFdey2nMFrtll/dauvGBZFys01Miihg+KiQCRSK6gmUze
EOsU7bU7TFeb5x0LiJ1HjloayactCYIDUimuavCZyatbm/QhNg9jXi8X3uye4b1MZqfNMMdAR6z/
UjSbgbSwLaWpT/KxzH7U/Ujp0tW4gu15K36OEyS/Liej6Qd0G1PCCt+zAeYQqRp5A4BS09yOTXbW
ypLwASloJPlLAyQwvEQBZBpZjbv8XRLRmQtdS++XtkjphjBvKVkfpafBjkMsfSa0Pv6EGc6Vqzu5
eG7mu7f3l2YvUTO9/F5kLn43kjBZ2H7OyYKYS9DduQFPrbJLTDDLkRRuSYwRfqmd+AZWjCkS8Q6V
g6E5X4l3JlRLQ3dxj8IsuL+mFk6BYD6Ql3Z5RR7N8bQKLrDrhKaXdwvVcYJj21ELF9qwpfKFaw5f
nMrHOHuV5fxkz38GWQx5TWVuDepHs3tpybnl9qz2mLvz7sEe7YYqS1UN7jo+Cp+I9u1ogAYu8W8E
gR+MTBQm6zxGw2ivBtiem0jwDphil9ggb82IsDJ+7ru21kXsFMGjR9zHLzBtja836/ojAMrYyVtM
pY2ztVfuVk01LmL81toPTGln1x3SGyQkCwCbT1U1m5hxlmgpvtn6/OIGsOsK5ffEFF1gw3qYIw/0
zIEqT2mxWoGk9IkwElQOZUtfMScLPtS1P/vCFVEitayrstQozqgdbWZFqoGYNYI8wCEjTkomD4o0
MZphBSxPQtrBEO+by+vioz/MnWLrNSEGqQFWLQoh9WSbkPbMc0deYiU9x/z/oFmStfLxaDk0qzNT
WVJBQxocpiwkkD5wUS2k28PAEln2SMnMzi8XC9gT8RaXh3l8Z3SKDl9y545GWdI+y2eG75lXW0h8
frTR8+WSkGcxE4IM7fEoQfbxQ4PuFqDhnQjdSPLMX3Zc7vJyUIR0+RSgPpTwWMaavKISVVmPty3P
sqyTDZywUEAXCB4jV7+eNwp9+CtIVRE0JAdCNzBKmV+edXGwkYFGRXhnOg9mMylEW/rMKK9ecFlx
UQRdFoR55yePnY0mZl8V7seska7a4qYcWpoyPFI6ZBLBhhwjG4BN1Vd19ox2iV3YXZO414yJP96b
oe3WdJTXsdE4E/i9kaNYDDsK4rNSxRKlaxXlYmZePo387CEAD0dbR2CPlH0HFf9ztSenu5psKeMC
vE4Na9XI5cDDlGJDEsxIKMJqZngSBtFpqIM7SC3CWiZbzw3i/6FJ8SgjfMe6CoagiNKAelZGJuaj
kYde4vn8jSaRv6FBYYmhW5lvJ5K//J9xzMU+ELEkZKPNI0972Na224hU4/4hx+QlSCW9TpB99KK7
UFcZMqkp7wCPcuUR6EiaWLgTlW35c1FhBXE3cToHg6gANQNTTSZKDjoDKJkTjszEMMPEbl8zMFbc
WQWSYueeTzaiKcNc2Z2ouAQ2rUtjiePw6ZN6HB9fxiUWIH425G8ekpAQXuvD3oAwaEr0Hikk7Mw8
gAMLuhdSKKsZt+dqtd5advSnsg/6i6R93X2ztomI1no7nM2z1HAPFVfJFM0K6I3mvu7+0M3cG3oa
DouY7StGo90anQp2Csqal7cKeJu/ThG/bW3Q4Duaatza9LokHmwr63jbSrtZODHYFbwgHGIwuQ96
/uj9EAsB8Tx6BWMkGlXw/Rc/DQ9GX5uF85RYUkubiF40/VEAHOQ3CluCIMcqJHVfK/TzpqYC4+Z9
fGZJdJGChGmB9VXZ3JpBw6//8NYKrxMVacme0vUxF7TTBB1UGj1vTl/afLuQ724MrIWGLHKE/Mek
M4IfkTQTXnnUMOhPteAHEzDb/28ztAcGkq9MIOtudkcsT4uzdYc7ZJ04Sp5SlDyMUgMCp2QnIS6P
ER59Wx6CqUuSPPX2koQG0XrmNFsElTGkedcrjd7PX7/aYlfaTT/922NOQjAAGvRTzVZ++U13OE2G
KAdNBJFhdjMpq4ieLh9Yjcr9ECCXbW/zVAOterJ0EIMZjvd5CmVQFCiNMf8sLcVkbYJBPSXXmUOA
FItRSUsT3rAkpcrJdeBjTPUGdzwfH83pfLpCPdQ7zaCDwzk0CdbxABZ+CLbpsf/UxvNFVrFgUb2q
1enGfY+HlVaSTf0v/YS78fZX42j+g9SYbCSUDsmNV1HYMqXcMkSCfjLrXt4bLz3HFZBhQICt92Qf
/yAPP5LfjoUogl18Lstv9MgIYeGEOhshdraerHTKVkQzA9raOOBXyKzkGgae4DOsAqNTkQD1mtBK
mIUxIlteWVxzBwLUqosWqjyVZAWlm72qzk+SF/dvDrIu9p55inBmmCXqzG3QGyhLGJvjfBbcRB1s
JC+MU4zw+tqtHW2j/lKcmyIeaRVB7uZapHUQALvakm3mwVt2giywJur1WQGHR8zXzHRZ2BgX2fmu
0mSAtLEkLZAAZUvgQg/Qt02qZsRmPgI3w+r4Hfj+w+Zg7ISN/1nb5BlIDE5HvfeQP+mdpEPmwtfR
Dqh8g2Un1U04TPmBXCq/hSQui3K0dYlG8zMdFePQ6JYhvvaLI6p0YUqVzLhAfnx+L0AeqxiLk/H6
MYu3uwWjOXALHiDHOB+zeFTB15aNsBMq7hPLRE6X2aXzhviWw3XcBTuciOWI1M1rjTJkE9+TqCK5
lJGlcJ4576q5MlLgr+Ivzrt2b4M/rn9fvhvrhniPaKq/8prf8XALFFnGNKmTeM1LRpLhp0JnwMM6
Cb3EzxXNJwlB38iB3GXFf6B/0ukfTtIo1FZovmCPxoyInFa5QcaVL/LHzIb/shBnTU+x0hZJ8PUo
Yrjrw2l+GJ84oa/s1mta4gcKdz4zcu6h0VnVEp3KkLM5xaGBams6RV8D3OGIO3rVZSjQ1aJNsUb8
l0S+k02yJAbUlA1euMx+zz1BysRcsPdImCnMzZTSnCFuu8eVcZuoNw+nqeYu9Abloy3ZfU02rZPg
BIV77G7tThSCAbQ0sh5P6mr+0/+N5nWuFfdZlCh96O01l1adA70pbFDx2v+C3QDAMzgCdiRGoX0t
bLm/48u6LsTHcwWQBFvG7TduOvBEGHpRYs46z9yP8gMN4dDMYWr0gLUk8pULVzGE07TDIhsdQTxf
E9QcaUeu3glqHoxacfkLHuERefSTmY0ewATzbOBMhYiYPstH5PieWPsxTQSUSjCN0VpRZOulXDhQ
HPMVNsszvpcZW29GAeNuw9TCe75sJWAtjqgy1ffP2ZeEJW3HZCWq2ZARaJGsnrqqN4xxRQLctKDP
oy1UActb5MsCSI0MSUH83B/MR0thWZV1mbZXigCXihgbylJg3asKIcRqURZbcdhX8eN8HohLHxUv
Zyfx6Efc9Ec6SYUQLsK9bDlDuNeOau2tdEv+ApjaL/LuYLyfkXp6xjoNG4JnbeZLWmM2dX7+MNpe
khT2WWhHzdRwrlgJ3TCXg19JtFUEFTT1PLDsVHbRr7Q+61ECuwrOA6jH4gP6eWXWw1a232cJpsVB
n0We8KitWziVRpJB3ll9Sp+97THM76/L9xFzi5QZbqAUKVZONcKtsnblQZcC+GC6cTPHdBiD+Koh
z+XGzjPQvWiK5dRsqcPrBwpdwIHuAp4fWrR0d46DLv7++/EZOwU9/+KGqp8FGek2wcDMzFIgbnHP
UebriCJDZkwiqttpu0LSUHE3Xc2SkQheUavNERzCQWvBnVLPORGuHG9NJ1i71xnxAaZRxGMY6S2G
ZxG34KsmqpU+Q2wugkr2T0nYnkvB7Q6pqQX86AWMl2kgatEsLqSy4OfaayD3+idyRCrp1K1csY3e
tkuOygpM8vH9BY1ricvvatuzE0eIb1e2CbghuwTzupVB3rS7mPmFq6IJMJN3bCVjCOFbo58BLiAG
zTVIdaBw9SZ6FnUZIXpXuFQ9bx6BA8uQU2JeEuHRv5clLb3TTq1/o7TH5eTW5opfZSOlud8JRvsE
uY9e3NZgAVRvZZ/jD3LxqaSgKgkPSn1rcZ2cOHIV1tTd0F3wzjirqR5La4Svq4x2rzDmK+aFCwW1
9Dxmo1GEoAmhr1y9avEus0Wqe9Sg0GlLEC/kxp9HNuOYeXqLx+vQKpFkkuYqDsr6ylbebJOQmc7K
j5szNd8zzrBooR3tojUP4nuq+BOsbAgsi8U94QFn4/36TcCKUiCOOKvXDWnOkdLqZOk8B6uk4VQw
g+G27H65nGqGmWoF/LUgxw2a4B0nb53e30qVA2tWD2b7KmnAD8DJeK2+0npW3aOMJyjB8GKsPhYe
O1SZLMjgz/V1CoKYwiF/1WArg+grmVU0PiPCmfhiAE7RpaK4HFQ+cJM6+da28dxceia4jNv8A3rN
wzZVApTDdCXlKMUKU8qZbQIYZCn4UdkQAa5iPylj1vf5KKAnDHWGPfBdOgqf5nqX6Vd5L0QcXOkw
HuPe7YFzPWvoUO0+2+n8b9GhcFd5XHi72G9w/iF4gM09G/qST9SCq9IufnbavKpUtUnPusb156JU
IYqoZOVwXL07SSDme1THE4/sHoO3bXtR746aI2BMMcPNAn9iEb4quSk7WA6/X70JxxqIwvEhv+TM
BZivp9MM3S8g10hWQC2OS2BTsr8Cn9bhetaPiO+4WXyGaMu2kiHrqFQP8QxDokX6J6v7L6c/Tqoh
uc+hjUedc3W5nft+WxhFydReUs+Zn/4NaDZvbIIYs6t6irPeZTXPDIA4/FXzlOGbjABDqRu9QKYk
Ga2VwK52gl4y72+92ztJU8xr0JYQgHOdAhKBbxg4wAah/rodWLDPX7MNLyTioyUJ9TF2wb66buN0
WXejAO9VMIObMBeyTB0vVrOoD0LwxgJqrZfdfbAh/BNtW2W/7xZohkM1dK810NfdX76pZUOlj+5T
AaxapENzNlHoguaIALwZmoHqE+lQovey/fGPIRhoZCtCy9HxWdQKJT+I5HWIjNOdBJ4pV9AeSLG/
hfIvDm5+TMC01tiIzSysw8IiwZfwqq0Y2AXIQ53IhiHoLEbwjipZF5cMVODwIdXzT7MwbInViBWq
b1N1XmCgk1rVXqqcin+eJ36QRFYWnyYrrl6eF47VU16c8c32u8Ufr6ve+H0VQ8J4hHnDyMS7Ov5S
5jtBiR9QOxSvIMmeKr0Xhb7p15JuEkwoGGBwO2M3K7cVvgHJptGlGCzyOSqxPmzW24NdwvrctjEX
+Wl8aH27cVTqm2LgGrImTpm5N/1ECB86r0vxOru3XdH7c8CAPl2GpAXSdLG2rjOiH/vPTTJdj/yA
AmIeyzTw7aZFKy1e5vKI/yVPbtX8gQCDd9jFWJJsQXBIm/LX/+NN7IWXOVd7uufKW8ciWapuLVjP
C/6m+x8VTogWrEmjeTY3klveCCfWk/AGz0QzzjZAoux5xfG9m9zWQbHhhZOvdasCoRIt0A1Jr1rx
wAbzsKV8tlSrjOmudkv+U6cvcAjTujSvvtcGNweQjujAxWFhn1o+yQk2XaOG4tuVS+QNHWCpqIAS
CD6l7wV90RBoFCvYV7GqA0TtcpijMsgSltY/4JTbQ8xjdBXPrciLPxZi+zvaSFCskz5ib2Uw7TNz
AkrvCTJSVWBcFCpTZVtRsVwnYocilFEna3a02ENNIV3zzi910VPIy6DrgndqJ0aNrDcYRG53GqQ4
1i2ClI6eOB5ryfD8MdgEv+1wcNEv/tMZ0kXkNJOco0ZLodu7+KjTwmPZ1sqI8EjgJT1i/955OsPa
TaC8fxVdGVMtVVziS5KZrq2FT+CqZc+xmT07r0Q1KIxWz8RnkOvvEi6aFvnHbpVvpEiVbE+qRg5x
uVUjXZR6ewReM8Q83FuqBUA9cc2tN251EyySg7pJyqqmjQNYpw2sl6gjpq+k1dB3+HV2P8H8ViuJ
arn4dm3OEzj1Y76ksV1VT+RDGZoGsWeBVZE+t7ISD+W7wkq8UqgWKrMTi2Wy3R/X6ShSGvRJK2FU
GwDBymaxGdBaD5FGtthi2rVEH//FcCdYRTp7fbIN6RHBBN5TzN6ENeG+iWZpppUu/KO5UVkcNJhf
zIUUJqvmYngPzKDcsCHZcXs3QuT8rO6VaHZ5SxApXbMH6I3ibTBv+O8xmK7wxwwUi/byJYA4GCX1
0/Jws0thu0Ab36tdBKcWMVQ5wFBLoxC0Jz/Ly1iaLPdhwCnVHLazuOcZqjAtyqBdnGwD7m/YORNA
uy8+vl5vMuKhezNzqQ/M39W2+qshg2Rh/X0lSImEPqRIaxU4ZednjOeNrKAQnBDVtva4GoYMJqUw
+cYEKXg/0LooQxHhh7iuJo/6OKQ1rLDzNKlynHDsJU/xy31Q4IAHnkOlpzAYgDr8nl/X4ypSbLYz
eNvUllAfmyhYJnRPFpyGeqU/YgCxOJ6YUDbLTY0QZGsOFa+5uU7QIXPk8DRUkp8tXMGhOilmZ0Di
+ZPEVfNw6t7q/x/ebQBLlBMin3XTf3RxtXksTUrqGCkW+9FBd0gH/rz7BVmuYbn+Tj4Ivtjmgp0o
vKCFiU/LKzCgcGLuou+VSMZ8curCoB2pM1feVoCqZt6GBIqcYy9fRdNnjFpRqq3sLfjrqF+XctQw
+73hpi0S1p1iEH2jHiUmcPk0XcCdk33IBiY+5VPLhQU9JKVlBdoHIsAIi+LC3ZTvDjpHMXGYqbfY
EbeUBBXeb4+HtK25yMY1Kbra8yIfKeYHvyjyQQYcHmB0C0sdyR9iR3CdI5i7pZPTyeiIlXQZZqIO
Wi62bnvvDkB3ttj2lacT0elF1hUkiz2umJUyLqtRLe9lGfCro30hMNiZSCsLEeXLl4joJQm4NR5w
exvLmpzBY5cu3tLSjR8EOnitciXiVctjKyqVnzzFVhqfRLIWUvEF7ar0BcNNC3CBohxwxDuGdktm
SCQqPhQ4ciS6m52xp9+kTKcCTGQrEqY/a0VOi8wJyFRunX+pdvLrAbkzFKd6Gm10sGHJ889Ggo/O
fBkr8IJWw7tN0JI2h2PU31Di0eY9IOrCiFkb7/Z+pj9oxsF07Tuiit5XtsH9rEppS7wt9rGRfnmX
+I2yRzuoZoh+nzNv37ZhPsHK3eigZNj5xLG2RvEj880G4xYgVFxXlSG71KiKqairMi+xT1bW/2o4
nB/60n/ycXBnvsRhR2wNs2SHx1W5DBIFGDPSykx/LLRaGHuFw1PE2TemXFLkVPDmxaNve+jRFcFz
m+lgCE6BhPqUZPwzErdU514dJFmpHCXnvCMEmzumEV7sw0FgAVU0BU/WJ9FYzUNwN+9yV7KBeRnr
CgHVY7RI2VBNqnDHbHAUdsjRsp9e+FXBgqDeDPH7lA4cFhOcsOGdzdrh3EhJEtsrqo9rBPnSsHzV
1SJ/FdjGZuj1XwDgB8tyQ8E0hUEHBcO2ozAC4WpAS2xIwOBOxvRLljAzSSnV5BO9NMfv1AOPuaz0
sjEe+fhGDDz9z3Yp8uJLfNcMb6/pdnP+UC1h86QiPmIQ0V2Y5h4EL4OGB89+G7io35SkNHdjyASo
cTCS/LkZ7EHUC0sZKCDtwhWZ9+viyfip+Ktl8MJdlp/Yxb25SEFP0t2cUKxdzOpE9eZY7VPvItRk
JWQidWLT130o4MRCf1f0ahW5q47ySJWg0Em8WHucK7P2PsDJJ4V1+bx3rBXR2LmteNsAZygrhXko
HpkuDWMUh5ou5BU/8XoAgCw7prR5/FbYltNIoEC37avMh7GXjLU1wGstzDjnZK5rx7NDeha3yZ1J
fPSDlC2YFY32DesYCgj56XTR6N0uBI++O4C8N0ekbNSxqVjD64P4YiQ3DsvjhaasJTZkn2ZuARYu
JXqivV+Ho4+s+yqlZ6yxn1Et9qJt1oHdXvy1Gm2+UnHSlHBuM5V9tA1tOEUY0V1nT0bhypvneX/z
sdwD2h8Si/wD5dmCDooifCP9+M1kBftCuz/pv0K4dBqNhnhd0FGRK9+YExtEuUTM1ilLoRNMxR/t
b9FEosnuQnbv4TEKax8oNlQhTwo9+/mTBF8LcrwFP6q18m+FjKdj+Q4SIdkJIpdVh6BVP1V/hDie
m9cVjEnHmPSHpb7EObmERK/e+F6AKr7sUlJZ5o67qv0Wn23zIVUOSkeheG1VaOu+ytG7/riQJNXc
R8kjPVmU5dCr1B5AoDgP+WryZ4VnUROOG12Bie8WYtXY3MUqLb9KRU8QM5gLhJFRHaQsSAkT/wDx
JrQkNMQcad+TXpWzBJ3mw63lvN5TTO3hX6Ixj/Iu+VdBkAA38XDdnffPxMQkKaxwBXPYhLgVp8+S
pTOIirJgqwlHKvaypiahk09Q6tOnjoGl6ZaoHGq1aGWvT2cIBH4T4yjkTzrNPjfh8ir2pa2WvsOo
qqKP4EpqzOxrLhH1XN87qrCgqCdJEIVAg2iGoAwqLB1EmtwP1jlqp2/CGoJTX74EQ+Mb88+dcidi
1PGF8ycb7okzYnH6jWgFC8QBZusnwaxuH9UzyKvnPBf08FguXn3KnOqGy9dfPykGsaQlexYFpoxQ
vvGrZQeq/t3DRx5znZmK3p95HlVtrTl5VuOPm82Oydk6Opl0aSY/d0N8GB4sDY0VHBpJhONN1ZVr
YpXLYC4x5UAedIlHLugai/6bIiDAAOIA23abreTEhUmVvSN4nPEfp3P+bLFTlRLCDnxDuMKa8F5b
vNDiTmtbNoP8M683HDjZ/XoqjinLkZw5CyEGPiZfCc7wMqya/C6SlC+XtQCMUu77UVjsJkohdLI6
7nMt/IvA/t0/dcbL6LH8BqGdd37j/wQyVl+qttTxgOQ3jVXVCTl1gFK24aR9tFNl6yTVcUw6Gswz
1lJgiweDRhoQL5n1earGhHJ/QNZIQ1j9vJHXU+7bbkokXykUutaiiGzS1SyXKuDRVctyCTARVNV5
+mntbMHvNMtI41rswibaaPqOSLOR6ThROK9HlNZrYKiYDFxeH1QgIIP/mNVnO8gGsfzPZ9THbITq
s8Ks5kszuPSt30Ub7xP/xRVLsGRCUXzL1vyqB7aH0Q/+H8A0jv4jhZNFjJb1fI/j7Dogmy3R+sHX
J9Oty0Lzepyfx/NBZ2ig9ooOALCspThGKHNYLNpfMLiIMcJCefpAMBMwU/Nxa9960XtrsY4N9Xo6
aHH5h/OiQ2Qibui57GrnNunbzT/CB8xQGFF0BRr2jlh2hHNPjPUOZdg1C477x4N55Cc1X77qSD7J
xiT3C1WPeAGPDoZv2j02Gfb6fPYNPeMSaGSMLz/sPXU75UFUyAyzSO0wRYDyjey6LyaxnaNDGu5T
vBpUZmhkQnHEmNMOA5jGWd8VCy7ZNa5OsWrknqTK3RW6YwH4CQSyPRr1TQm+xkxyfPQYdXeYMlPL
1Zz2MIjtNaX3uSaP+zk7dO68+kt566r/1SG40WkpSH5klyotVPd7eE6tJG5+XjK6MFDLYCbFVIOt
L9kDEgby4MfMxpYvgM51UjHqy0avgnMUefReVk7tgAm2cXUi1PPrWWxnmQXy3xStnK1vkDKnRlRu
7SUzhh+FW00ZxtP3odBIAItIGxJJtvW7K7A3axKWXJa497MntxpT0iWdFCSINqKa851/+XUFOLYr
sZ3gkfkLrL5MLe7W8XiWVnPHxSZV0foMHWRVtXQ6g5i9qKm5bA1pNwdZtvKUQ//vGb+MMK1aY3Rj
OBrtbmd52Cy5QMM8XO8lKBW25jlRZS/Rqd0PLnv4s+RMku2ttDjhf1Je1SuOddwAmxUH4KSI6BfC
einE6eMNQpJJ2bv/eGFu/Eo1QGBMGVCBZJTbDJH7xcBMqMXmgC6vbxjjRMcFd4QqxQYCFd2kXaMM
NZAVBDWbDLiseBmuMPhB03DWkd/12ArHRnKRIu3focfH2uJEvL9tRENUDAyVSCfmkHdc2KaRzgvZ
SOyVHCwLVKpzyqJoetC3JKjtdgcLM2G1lC7iJ2DKxln7QXtuVEje8XmbYotaRBtXwr0Hg0Nv4AOB
1dmLNJTNtDkt+5Hn296Erg8v3/y5skPuMQnDdij7jdEPnZgLsO04g/321qDO5G40L3ncsleQhxKT
oHW54wEKt3ry7zzQK/z+Od6IPOvaG07jrnypkKmB1T9juKe05O/c9DT6LdUvU8Uxc6+aUONj2ucI
5nMVLIrOCUl4i79JMpQhnNiSQiHySnq7J4NZrchGtsjsTwEA+ptXw1azqaOt/dG4z7pfQQdUVNTQ
qcR4b5ZJt66SyCj0ctheJTS2QkfF+GNK1IDSey0QgZUxlMN88WETaiFEOXb10gIOCr8vF6xjTryL
8P9rFiCEUPBy93Wp8kKluKf/MDu6y1SnjuVQYpd6XXgYa0iag77E/8xDYHt1Klo3mOo35Rb3TyqV
jZMjC6yWd9yPIsnbqjKucspCcpmn4Hk8BCl730sawRIA8MgWriit2su8cpNZt7TAv7Ji4mE45ZuH
h3WBhVUBWaC/RIsKJuxazGOSctFBq10rRNSvlfqvX0ky6gqMfXjbtGYOoKoohHedUhP+b6i2vgs3
i7TYMaGtIaolKQPr7tq37pXqRgTaxSDd2HIAq8ryd1ZQ6RSntEVoNVsM9jWJQbz1uZNOpOlRghtg
xTSPcsA89pRZy1FgL0tV3DkH3vO2kt+e+gkeByl3UE+raw3ePVQPU8tmK+hWaVxNZaOMx5qHBrzl
0Mjm6wwQSltlka+9mVlDJwkjx6DBFB54tIwDedw/NZVSP+MEtt4P5na/eXt29/2NyxFzfAzt7DRH
qgupkF10uG1s8V2I5Wr3/fOt1FskfUkYwZbhLBWCPbW2vfzAtJcuI9oEcewKCGz0GzPiab8HtwLp
ITm8Nj0a8RVXNhfSDr1J5kIYpviDPKfY8kFQtSdJ3JBh4FhmVuQI1dojr72kNJefnx7qz80NEWMV
1vCR6Cd11NizWbetfBxNoh/iGhylILIht3xrs8nXWxzm4VKkeofA3Bp9tA0Xusn5oYUmewf83Rvu
Xit5wTKiMMefUBj2z9SWeD2wplZaBFEjBUGtsOFdfjAM93JYYLRCTVd+tje8lj/TTlbNhLM0Kizv
9Gnv9Ktvq80/D6P89DHSiVDUdtWZMDETGXbNJCrzQti+LzMq0M0XPmSikcze0zDd/iXIfINV+7/G
G0cy8gV5EaQNRcpQ96P901Hksadw0yFI0e9s57Tf8wWZgAwNN0950GCT0Lt2/LT8hKT45n2JeR1j
FMD0zdo+zW63XtC2sna5q5MG7mL4BbHx+7Ps8NPREy371TAa+t1egQ9ehdyAg26M0eqV2rW50AW1
ZSZsPBC4BAh502nw7tVUIRfDRSrxgKBKkieQjdZBbqGAE8fydeBLsLnOmN5lI1tf0Rdd91/s2OnR
+lC3hww/Io+okWSOfEFqDODTeAyn3cEuekZbP3LjNSsPd8Oa8UNIQkfoUEBet82axhXWeIPfMK1m
ahG4fz3Vn4XYAg9Lkon4tKWcFCGfBcLSpXdv7x+zG13/FCYnth/bgCq4qU5R77+i1eNoFDJIuZ6E
WBq74ZQGyss4lnsaFn8WMXGac48m7HaRQLqKlDMx75aOrOZHHqyJl/xelEsTI+lTwNcSo21ELH2U
W5jAv9hIomTxaB/3UXbk24RySoEyd8GQuZmv1X/Ap+Qb7iYWYNc+sQwWzvrMiiR3FnPRqcJh+2vS
i2bDriF6nBh0vnPakWQMwtnLKTJb5PuBEmaKo1yqu0grT9y5vGc3HBXItiXU++bhc5pf4NS2bvwY
3U0SmEqBUznZ2vrj32talUlYkRtd4pYv8AQ3CPzHCg1EyiZeJm/AaCVp4bACqURl5heuNYY/l0mq
0szUNxbB1gB9F5JULo3OpxrMNmkq08xWUJffTEcKvgHs6ximuYN+YKc67z9GOs7deOgZ3+jTe/QK
YcFPqumKsK97OQpOtttp+P9YQSwCoYd8mSofKubMjV/m/YkI1XbcvugbyLxQpKje4Ay0WT5kySRI
m+NmX8Gjx8u7snfd6iXs3LQO5TSlbaK+ZZDL47hMfcMnR2nA+f0FrTq2O6fDQMoU2YoLdwus/x7G
KiyNbRYqdjY8znIGYKhl/qA0X5GSFuIghMF7xcutuva/8UDzH07MqZUrSJ3TdOry7KGzxv2NGv9p
vmaePOv/O9W3CyW4FAZSQAUl0zdnHL7u9BJYMZrA5cbOitsphl0jwE0FXpqe7BjUYjyMxSEsb4pD
268+TTVKblBjUK/j5SXEg4+36Ymb/8CxVVjmAjl+R+od5QgIs7nf+6Pm5VbjPKjuU8Ev750MwjfT
Co+PZqZzgji6nI8rTn/NNgt/GEfrW00K2AsIbhFw5SItR7w5jNJ2C8jgzN8p1ajP6s//9sYEkJ7p
ZPhcbNRUJGJDIXSYAkazGnzX7XFPeTpmsHneGoBU0wTMsn5gTvwahs5vmsAGzLABreVyjAiffVm0
wsamEokbiLhplwUju9QE9qWkduBQFobsm/s+SX7xLy2PZd0mVQyMkg7wmv8+yrOWH5Nlu6tM5ZCJ
5VUcOXuQW3xsT/s5a0alpazJGJ/5dsexY6u1/JQ9KX1AVuk9XYun1DpwSueoEXcv+SwYpVrF1+h/
Gm0C5m+UKZO71lMIIXP98OZTgmBt7vBiox7IC06zS3GCo3tqtU7QiJNP0oqhybu10kP78YnofRVu
dURSkzjI2cZTB7Ee+okPSWH+qV31AKVVZdeptFNhvHGWWJjZ0kwnBCEDysyxLlc3CEmHd7BWuivq
7sFm64KJib5a3wTtkDbu+E6Yr3Q0JhPowyk9v0JOqWIlB3gVedyWHHPPQ7UVkKoV6AMfsST9p9ye
geqwRfggl5yVgZsZsxmN+LmAi1HXvqhuKZJiljXleDOV8PZJ6//Py7/Uoy+Zp7lLTZ7+HG3fIwKN
1pXgjnFvpxZl0MrvwVDntE3e5SWCeou9urWL91u9+AYYAn7er0QGmY6M1bADKgWMvcpsOcd/O43C
vHMRGLIScoOXsqVfhIz5ln2AI8zJO9B39Eh8E0bNrcVInH+Uvlzr7qYdamYsrTyk6bEAmTQSa+TL
87vd0U9Q/yCXFyfWqAt2BNGviO2eJz71iWSzqVeKfPwkpFT2AqgvsAAydjIoz9q2Zp9MVdOKr1wb
diCcb6l9DZV9dEA2miuLd3q6wPDC2KUGULPTxA2NjxaE9O4jkoermtYvImlzpizVNQ9bjkJ30GGL
DjrUXA8Jqrac8+uWpilBuLbob4dV6lBdfwuXa7D5YrNm6XP2i56TsbVBvNPQyEdXRchRhdwVKYOd
lhBzBndKncoH+GTPW5fMxvs6APWOOYH7tchz42yaRqaL28nCAaAHmPfx6hT5ff5kW0igrPAopOK2
euhRzy4at4H6w+xCmi4N1PtBWlKz7C48RjLNBUbYKXJsY0EC2fIQHqHoMCQbJuQw2ygNV6m3JbQM
LOlkZYQL2FD3uhVABdFAUr1NwFB6wSFZzfLSp/CWHzTi4k9mDDFwjrwdCmwV7Z24uYISaT8GGEWK
0jtPgVxi1VAIPtcaBKBYSIyCgykcRq7qRZbxc4HHX/1JPtCs5SLKqOmhZlW2x3bo9ehHB6Kex+lZ
dtqn1426TqZNQt/mqAigMLXm0ZoeKn423eHfKLh+cFp7DUhnwabT4pEomZYu55J4g9uBrk+jLV/I
P3/tQJE+UrJuI8msBGC4q7jlHnMpAVaxZzK5NtKAP5ahAzHVbtWMPA4MbyE8soIJk8Dp54tey1Gb
OsSm5WxxShgTM3iVFtXRb984VI09/1Ohnl/vvgUG8aK4+3e2D5WBCT3aKqhb4s+KPaW9q+RYO3+R
4khdMw6KNkkYqTl34TsvfLonr1WZ3ahFtNvLTHxsoVtMDsCB1Qxet72oosBqigKZnWqhnUJYxSq6
Xqsnqfq3MNaiIONuCnMZnJSVl6X5Y+rSvds9Aczc9SkN1zGshLi9eqJ+i5o4/bJuy9/+57RK42eW
iRboVSRnCz/Op0lY+M+nYiMve32kZcxnV0t4Wkg44T855S2K0jTDBB8yyA6OP/nk71U6OZ/2KUCR
ugGIfmAj06wwfDrCnXbXpILZFJdDnq15eeTy3zdma+SHjsDSeutSKJZaz6YbkyjVuGivJDt2iYlY
Kt8uCnEyHylDE7N8IDwYvUg6nawkiB4+xWu/jJjchx8gaal1l7jgtJx6D1tfEEd9TWAQ/UEaA+4h
BiV+GIwp1dVVtdr7hinKSqwIy84grhzaNmWWrewLrM7YAiXHGRw0TUw2DlfOVLqHP/63rUo6TCli
XaMq+BML9Rw6+sKHOxGPyWRLkFREr7f7DVmxKpl7+9kWVORDtjNFIn2/WuC0vQOUv3DvhVGei1e/
L4w5y5kVTucrOOL5qSMKgRQwSD7u1bEGfCGBDU6lu2jKF4KB9iLNgF8FRDuwUjASGyJ3P2x/QHeK
EHZvq/RApaq8BOTNZH3b/uImxhO/jgH5uBwmV5VKtu6ChoGIsWSzbQeuJDlervONGOChTXxmUg4n
qcjqOwD/MuftZEr8W++AKSmF0IH+/3Dak8nCp1SFqccjvi0M7hpJPGB9dw1L1sFulArqH97C030E
5Gdw5KFqfc3Qsy+9ZB2WpqwO99SuN9H3N4qzuHwaS+0XEhNLbpaBnNFd9WjtlplgCd++m+HFnTql
WhMIkynCt6Op0szMaf29+ACYjPl+AwU8owDF0llYjTV204pPEAhyM8pOPyUCYl0fE1R6BuK5MlX9
1/9BOrxKE/Bg+8t9Va/yTIyY9cM18Lj/NMLthyJQiPfzX7sJlIqj9sn3ilEOhTRPmLEp7TW3OVpw
HPqQeRoDc3B92vU2iYaBE8jz8nJOFvGGmMhuIuO937wnQnNbCeOwYOrU8IedQL13XZ8vXjuvyLXj
C50lbSVwdiCK+gnpJNSBuM8Xxb5gg2mikiWcWY3/GMfXjBAJNh7tBvEpp4BiF2EHmAg6UxBYO/O8
57VZsKb2aVq3V/UoyeHPlyNPNVV99vU5s8Uswxx7uD8rqTa8rYejLQrM7Bn9lX/jgG2fnIqTaleP
mZ7bPblIt7rGD+rwF8u/4kOSORj8Nx++DrliKtfZiSXXs2oADv9arxBWzLjuavKeRcvrDAaB0Zmo
UyoVQNlmEtNBTXtgg1HbYNQ+8P8761noV1GBbysuJLtUPmYzj4iS67qsGwtvxeDUQh3/j/aurYIw
6Aui//XuYWuMJf4pJ6+j5TEP9D9iGQ1TzE1uhKbXn4YaQgEHT1C4m0DM0nw9d1Z77QMFmjcrGPvC
ngkuO/5h0L6ELPBZY25x+5W6yI3Ok/JkasgQ6Vk6/9pRKbxnfxLJy2NWOpP2sX/UhgxS9z8cRsOu
yeEaQeIxCf33fq300jlgUeHezzpdjq9gY4xWznmdoYNWSFDu5Da3NTCpk9fVRkgtNILpzMTdU/QD
LooXXke1S65cDBE3YZStBdVr4Knkax0P8sOmdyBhUiXWVI8a2/6Lf9l8FDzJym2QOGWKo6Vn3XDR
vTqAtnJyIeBlPVq79E3Y62tGZLP2RpJZQ07ZPhEB9vM71F6repDodxbyEUvhOSVVl5KK79wKB0MB
Kamn87CvZRaMCHXDj1ZJ9htOnu9HSD/2WKi8obLRwtUW8uAg+vxGZRDnSIS8REhcWSJlhfd/Or8q
lhCr+N1lelan7AGm2M8pEPWE0uSGV6KZoeg4/QzJwYBeGDIPO5lSxj0a7CvZYxcGaa+zCV3qnwNn
wyjz0vLjMZkNjm83IPd0VO7CsXru+jTK5DFDZAj8BlCWcPEijEeKzw0sF5axEZ/sDt5iOtVCf0kR
0IE1wIsCESN2w7fUJKnIsKuf1lwpd51etYazHGHudf65u+KlHprd9e2bnUdSJyrUCSu48I8yjagE
sGjt2eVXNxTSbGiph+9drDv6cn91zIRqnPuADAJNmDxCISvdh45XH2Im2WU56J3cp8AYXWxhpbj8
5QnafCHYQq6nhDYmBCzwA9BurywYMHZ6pxvbCNvCYj1VYg8e+kp9LMSpZIOwjPFbsor1U/Xr09Vv
E/VD/ch2Je5S71aDHZ4KkBZDoi0ikNX7TovAsI5zaxtR+v/LjfRVr2eUJW8pRACRRlK7SZbMdVNy
3Of7km71DCA1fqjhiYVChdhTB2/lhRi5nIKOUYFQV7WJIbXsHvdSFOzDvTLwxJDlPcUzbqiO/S1I
JkAP9F4G8Whr43MZVznWics/95gYsj3JQoTXgCiPKcHHkk9Ctjx54AmNih5yQhM1JgAX83vV/CQC
3AjoCW3q/BlI0ryiGWCxqnLQbvGqrpYA8YhF3xY0mjozGqt3L0wCTHnklKAYnmCTc+VXMtwUr9Gm
XPD+pcHu6/FfyJ6o13tIoUIQjmLD+8CcVoTVhwKmAfpsc8wSZsJTPu6KAdo6alyz5bRtkWWsXslg
WWCTnA5IYOwMMXaXt/ZcNdht0yOyrTlwKJTChoVXb17HbB1wGPXjF0UabIMHZasxPV6ddPbhWMHN
POR8kedOulBSv3r02D1le32t65+rzggK5PTMaRnrbBn1oD8M3wkEvfAsnDYSlIiUyyf/bf471JB3
Sby4054l89h6Ii6c5FfJYmLK/2YEsHhzUNEGN3YRkOJV4jLSt6R8q2hNt1/8t8CgTwCSYupcJ0M1
ARyfyKLjf6ZpcGWWSl7rhPlNYlLA3h6vgbDAstmw2VLxCsxHDCVrsjAKoLhJK0GdfOAk9FZtb7/K
qp8+ZXm6wrMm0lKSilUcHlHDZ9OxeClyhn88XsYNvRpGi5eUGR2iZytgx8xFXsyP8JHxg4JLn+IN
GJOL/9cRJPnPIbtEGX2r25AXpbliqy5qyEkv+hZ2VsZTw4vSwPLpLVhS/fcaWi7wi5xPhUSNTQQT
6eSshMgIw+aIx4ewxG4qQy7ScA9cAvFqHoJZ61Pn++SyP+NuqJgY2xsjmFMwa1haXaardqWbcjY4
KAMsp5XSsQZrKg+ks30FoD/z4Mm+uBMdrwq59RCVGpHwiXLjxB0TeV2kko1yX+CztnwpqLuQP9zd
Zv7e7IKD6wAYuuNzmvdPxWy2rNr1KRaNNdBtbsHi+6rEu+WW46t5fN0iG7jaQxg54MssHJ4Ch+2F
d6TRzS5yCO+YnPEQezjdiNyq1xyP1cPydx3ZsgRjE0d0lLjCo+Flbm8LReGmaHOGX4HlmWktql2k
0H+fG97UAtJaOD6iRkwKrqmyiqYydu+ivYPzHIRGfQrBwuSCylk1AIzcRalvSZjMM/MzXVHdHxH9
83PxXjE4h6z8irXqcC3Hdi310p30oRu2AAKB9AN//EdExzSW9NJjEsreyGney4a0x1TTeS9aIvkX
chzul5uBh+jzYl/e4suAFttGEBeyx1yziIxAY/UbwJaLNq8nc7Z++QaFp7hJWbWEJidWU2YXM/xV
TpvyO6um/OA2jLiCJjhNfLwgyxp+PXOH8HDdLEkqCT1gzxhpZL1hiVnISoTc8ybjGF49SNRftFUZ
EVF9x2gi7xBH9U5WCYwITAnfYhAWnJq+w0WokilqccKhf7/eJs+ctbLYh7OqXnFBUVRPGK7IDC3d
ah8eHZisFbjkWGYjAgZVy+SulB3/ietGU7PeeDT08+lUdhMHXdllIEwtzzliqTbZJ7+2KVNpVAs/
wUTdUYIcfGevzrFDQHLNFFoAPz879helNlmg59Pu9uN1oTcwbf/Q1b6puvXJvDCAy7ngFRw3pq+G
2xXzFr+bWmiUK7RdqHWoBKAZOuz4gEv2NIbOyDgQd49NbG+xX6jwP25kXF6JO+9UjNbrbxDcjyvw
ovB/Ztx6W9G0xixR6FlA4+XYous5CiPgPP0Ca8CH0gvbHg+/de92EgM/nXmEzfI6jgAKt4leonmz
7ZK8Kth8DZ85th0F5ibb7fvXHUCEI9o5J9AQ2D1YA/W/hGSWAd9rNZpXPYH40xRrnJBszBvY6S9P
X1Ltilg24PQNb4+VXHYM9QOycpqqIOeN3LPQvh/40Xkc7F5xCFf9v0A7j+moEiAayfb/K4AG22UC
HvyN2qlfgAMubGTwjOB/HY2gUhCCYJLA3xuQNr3BbiGMLvdDhsVHci4+iGTj/uiwzszjBbkQRM7p
VsPni4ioCa7VHBRcr8MRys1hmN243vqdHiqy5tsxkG60zr9XgtIu434djtyAppd1pJz/z90Ieish
qzAyJR3JKOfaq1iOo8wVGjpN4KH7bJwfTHxPSqdQM4eCiSJyTrHJDTGDEGZOk7bSe9ivI910tZrn
FFXrWA85egywl4+2kigZoaZXvL/E0baLsSy9tjFQBJ2xtmO0fsDx01vt6gNMkUIjBO+AadkZZ+Rf
DpV2S+yw8+YsUIYl+98lfODKGRnltG1UwNj1HvIErBZnOzsmQNORwpelcX/4YhPqketooll6zDJA
EUbKJNFMPhgqUFvWT4NZ51RP6SlbsmbdWWw8LK7Q1HNvhdqWP8DENyGnOWQI7rBJ1M5zgPQRGA7d
O+Mka+630EIBZuhIGWlQNobbPu8+RD5hwI2wseynkV71Xsm2nv64gRRJyl+WnRTOezo1efBKXcFh
trXtS85MQ07HxzTnyK2KKt5t8TvnAdk7tvL1piFLTuek4DfdfxTvK5SBzmlkxgnZ5OTzDOAZSERx
iK1PAdg7b7JlQ0OePdjgpjFFVgJNYD7umKaZov22jrYSo/akkt6bVjWQYYh0KbUOKcZFAi1BmMOz
EI5S41ZeMnOa4+gDM+WMdtIRRqcep9lQBjd/KqmQ6C/VXSooGvd3cjeb0Ks8tQZ35EjLTmyPmle2
h1ZMlWqUNTGX2Guak8YNZC+RJPX22rfW7MS66oJ5wCAZENZJQMrPce2R3Z0YluJ3eRnIR3XyQDzG
XTw3Z/AwgqOppEnrJX+2E/aA8ydq4M9bu5YxTKLM/w6HJiLjr7wZ0Lb/jm03JY0T3n8RqNg3mb3D
BPdqDO7K57FebPavlzOMcWx8acA/vtPxo/DQSgZ/xa5bL56FmkjWyo4+fJvkmlJvI6ALVylpEWdf
0K0TOQm4eCzZesw0mUQSOiyKDEt8sSHk6eg7IY3736U4G6yehC9fAKqcPsIrBuldMzUMvuGBkmJu
0qt3Bf8slWk8woFdU6h+VCrzWf9RKleOihOYuQ//DjcX535qSRbGCZGsKbL4TSsY89haPMjUkW7J
Hj2EatGfEQd7+3SrTNWdwrdXeSPcsmBFDVrCxet4AcnVzZ44auhwVLR4fndxtMdYYWzOn8MDDT06
nx3UHi1WhnMzprFSnH+AWJZdPMF7maPc8g9dExx1R11uaTIvERtSeMklWOZm4tec6kun/ma0k5Wt
t3vROtVBNAa4TJo58TI2mBY1JFvjn7QftxTETDX29rsv/pfUuKGehdJzGqvGjKbcuSXaZ5N72L20
oKEV58495qB1tPBAMGvB/iDFtrVc/nya7rAsRljQ4MNY6+o7MabYBNWu6hbB45JexuVctOMF5kBB
OseQ3ZWn4zugh9GOFE74GvuNkwp9XHL+MZXM//FgBaHJxHI8GxmhnMP3F74ffHMItBrxUE4Mp9qQ
TfHT7nsNopLHZ4vcZg/Ail4BfiX2LrHaPUNSEXi1KJNmVfc6/UztJpyZaAkzA+qoSh1T5Y07H0/t
64oRGwuYYM1f9Y8hTa4A/XT9HsaGKMk3AkMc2b6/CV6GdJDzbf0o6m9w2rPlrUUo2lEbTEHwNlCT
IoobZrE5Q0ysaz2PsjjE8rmPH4M1+K2vho+dRTMyHBwNDNFB+fqRzfet7Xb9ZaZnPW/HAcqPdI+K
fUKLy+WzCGcfVw3FXHV1Ykfxq06ugBVKRGxH/ZQrY+ym91XAI0tVPbQdwUKoXanvv8tIFDC9XtgR
1oIk76Nzlyy1G9K9uyKd23rix5m954p9g4PCd6+G/c7lwR2lT12WkodbODfOxeTBWDYXcnYtMbul
g+hJY/z76gi90HZSxSO2in5uuLonigcCdvHU9l2NszJpi+X4NKBYuIofPL8B45aiH6z0i0iFbwtR
w9rZylnn8xS+VPt+buLldJYjBiVRaMxN2Mnyf+9dk6WCL1d8rqihBv7Eg+jOlyuQzg6TOiRoVBkx
lFQo7MB3dU8htx1NFJoVffo+g2vAH30opGckTq2KB4L2/I+njs63M8k1nKGjirNji+JtKeBAmGuX
Qho7x2RLPvJwV+uCMiM6UIS1+bRlx/JaZJ9WpzRSVLvsp5VvW8RxjlTU2ANyCGh3WWogeMSR+Iye
H1gcuJFDeZ8AXcZm2ry/EbkMBWgADM3/sCgCQ6P3esq71YOR5Gnv+V+i+LxjOpcnKyZgxeFxv2NS
uc2VTgR8N0OFa4zKSqN1ajZPS145/fbuzczzLS3Y/r/xm7axbZMMqQfKkSzSfFWrLfqEyG87Bfa5
OKQuJCjvBOTOCNr5VEdj1vBQRGg2YI1PPpCMiAhHA+YBR6wM3X1ALivS1w16KeXgawPIxWFwYp/S
/CigJ8/JvJcvI5lSt9fwihz4JVzsLBSIuzvkJkLVY8IoEBSCz0R6Fj8hBd8MmHpzZXCl3xNB1ZF3
zUyXlzix3dqQzRZF2UJG8vOLAL6deUFQQ0iuZgAK+emde/qZ86UMmYNM36EmEx8wK9+ZnAV2lf04
aAZUoEUl68lzjues5gQ5MwX0CjK37GT0TAVwTqU7Ghbgwy0oURwdqVGWzE7uwwGoOWwUdNx22hjo
/ftnTVFRFmq3GYV7WuARsF3X2iyY2oiJyKwGcDuwFaExqtwBJ4eS+Y/Vx4Kcl7jf5qwAMeWWGA/T
C/aA6sOrmHixcE5T4EB8ihTvbGtZGTQ4guwLa6QHl5um8cgE8vD2dInqybg6sQ2BAp7tJKLGR8D7
LlcKcWWevob0dQAzCn+Ok3doCgYFm3LaBhrJ3PwpZ18/i0cM0nHz45vZ1DqicDHUbTGNWsLvfs/B
GrPi1mHqjlqCpcauukiYz6l524OReXTpSxizYKomcusaqf76lEGWpRA6ZI8tSPrw8MDMn8FF7FDA
dMPe3hTjsin4LSghCaEgoYj2geLqt8Cayj1v8CET+nV08QvByhka7zeSS0bcDH/eGXAkfYSuMEfT
RVLTk2qqi6044H2T+WnZMePYZb/ZQ5gd2zBI6DLe6yD5OtGrEd0a2QCAzSBigEwHCHkthOalMidv
jMOnT628tpLNDnYK48xsuubFr6SSY1SxO000iU4j+1ySyxQFdRJjmE6raK5qZ7iYUaSM5TI1qZRl
Z0vqR43qKbDQk2jnEyz8l/8rtbe+1At9W/eFsgbug+atTc7jcRDe3R+I+2zWnnxBa6fQVMm9AGQj
czotKyjGqOB84gL6NbYde4OSKRuZi64Hpee5M5TWzHKgt9co98RzCEDsiDGqm2YpAK/HiVbqnwiY
3Zqai87gKWWTSCRhnDYgcmWSLCAZtW5u6oO6nmJmw1iWYr+PMGzdI58Ae+y8+FBjKT4u6yMcXXg8
qoHF4twEAtVU5dTuwZJj4k45vbicG7wrllGgBRLFS4uFoU3dyz6f6xCLGhq5qvPtATVSKseBX/w0
Oh4lRLhN4IRaZiqqgPj6/nSRkZBAC7nPIX748XUzGLrTUUMkyGOcH0kB4qv6ma7XmJfV5NgfR9eT
MxxYYjiHhyKjfXvr0sVeUHSGdAfmEf5KuqvcEmMXJMzZlZEUdTnXaDVBJtzw9URJWvh1iwBTzLHT
Qdl11sHesNjSUR3LiZ5Ptoku+3veEkQmYvtZguBILCO5Pxdd/uiKAJW5FnkP6JQ+EPrulbYUYCI1
DE/BwQlDYXj36+2q4/DsPCStNJ0Ft4fYZVvjq1ws4iiggZRkpLgCKFC6KFR0H9No9PwLDKCssT1C
kD1NwNeqkiYz2ljvz7SOo/USQZxaDgYUIJoI6XfjKMhcO2VHDajeKn3FLINQ82doScvAQ9nkf420
6NHPYTkcgm7M1QJ8uMF6KHl8WcGNB2QSSD+HdE8LSJhIaPkZv8rsGHdZd/+M2WVro0xtpKYioqah
ijOSgHrBUh4u8ZuVHsG4YDCM6SG5SNvM+CvV6owLd1twdPKk5LdwPSusX3waLN4VMIXGao2QsACo
HNG1d2G585CyrY+y/LPL2PoatdNvQTmZrXIVXHBkzDDhKrIFuJTeUpGiRic8fHM0ybOiXlPZNAVJ
Jh4OS31YN3k7mTycwwzNXUiwPlZ3nCz4Pm8g/pK9zaxs2nlG2FHyM7J5b8bL2wyLV2HW4VNrUmp0
ckmP+hcqdsZITe09tONhHBSPr0kDUntQqO7O/Ls6oy82LKevbAHn8xuwEnZH40m9Sb7FbxsTGOVS
VeHf+tY9FzFOIclCeumoi/YGDSwIpgw6zT3HqzQB/Di07BG77s+1MQs0kUEBY80He+wSoHdKtF3R
p9TkWnRPi90XlD6J4jBkDGByjB4QNidGSa1f+LS+vShyPI+bHahjiqoUXmfCWX8lYeDccpGE+T0y
D0E0zw2bEuqhlBtU+acCl0JYhnA7J78ouu+BfRd2qHit9n44HvTTADnnq6bc86kVH7xSK/atlyN3
Yb8ZXVagX8wWcgcPPUBZbYXjRGzV1qcfP1LK1u+YRLA2OHnklUfGOwRYqrwlGvhBMagIrqx8KKOr
vhl7jgJ/xo/PLPMA2NxuUKJN106Shr7bwmMqFzf7lQt1WTNF5l+LFPgHphHkkYBH1hDGISR09O7R
pJt/rkESMkq4sr09rOz+iSr0rCZQ/PeQPtlEqrV/Vgn13wYy4HspPanqhexWh2oGJ+FJFf+pfzFC
2ee0nx6jZHOSXrM5K9ff99UB3PxKc4r1ELGKI848jSF25//iKN4WMsbwXp/sbkLB15O1Gw4scoMO
CQdnJXFs1S6+gv661XjnIJ5PAUne57qaClG36QHaK0BKLED0yZoQwevmfQ4im9oL2wIfO81nRejv
cMpN+gFax+t0LTkhlgrShto1lyHcv/dNl1Ew0lCHRm0cHsuuek1Z9rvdk7XJ4EsW27qe8ojRPjHu
SCyo7g1dOhltnawsNfBhj0nAAd9OcvZkrYyTk+gCOf0BjEBNVKYOHPvD6JX5MMMBy4tSg/dKCqa/
rdWsnk3N6o/oV83g9GnqKCMvvQOBdahhgmqG83tZTqfxJ4vlofTZ0zWyiWFk3voFSWeyM7bGzcKv
a/LhilTQ5wCKv7gPGaPYy7qMJecqezsNGB+pKytj+eShR/vNnP18qgxSv2bcCZv5rgNotcCnZZys
iGmYeWUZoWLoY6fAw77WGbnN9hZzNvFKFLUxj4u10wkEq4XdM/kdlKuvZ+UMYkuntv8mDr9Xucpf
zTg26e9qP8VsKKryXoLsYpKgcje0pH7MKdTv16wAgXao60ItuT9dKqCd81JNC16ubHJRyol4quHn
+D0fKkvTUw9Rq912ZEIwlDtzQPFqiCz4hn3EdQ8rzfK4VL1JvhGyzJ2upbkArwpsDRJNVWA5EHIk
G+d9n3m5Bypm/crrl79Pf0yKmcoWVn261278pgJ+k2voBYU9A9fWKSpUzxzxbmyUmbKeNLDhOZH8
CVH9aMVuGwFFHl3Q4YHmTnrqsaV0EBHUR9B/cBAH+llGeL+llS7CNPS+6vPoQt73T/RCf5daKXg5
1HlYQKEzryMExj69/5vS18VjFcFoXOJ8cNKYXt0X6vgWc5892d1O3EdZHBcJ5HLJFBbkXJKa/B37
XeMtDvtDLy9qkO5ujUHfPQLQiRd2JtYbsyhFbVixvHYI47LvbsYwJi7lZp824+EruCGjHO4eehUX
DIJeZHEj6DBwAa9q1oxT1g9pYMufiTCTKIZWhGuEsDI0wuv6ejD/PaNDREO6zyAFZCuWF0GfP06y
PUGSj9jHF0S6GE2z6WAHfgjJlEdLknoc0Te7cc/uPYkOzYvulMAf/PDI3b0cDpcAnDAn+TpNXJPC
XXSL+PisF+ZGHVlhFhVrob4XNfcAFPjZ1dSVti6eA0hdDupeAt3zLL4SCfZ0YZ/2AP/cFa0rRbs1
p9+gmlY3KpB6l6DNRm471MdSeTRjVdXopVFN9Qoz8BRvuLTSM7wpdpRYqdV66z489Dcdl+VAJv5/
+076vf0SYdknCUgf35+QpRN8O6Ax0Yk/JRwOxy9w/2lyeg4BeJ99K5/0NtBu9UlSZGhJ8V4CT+ln
K++5JVHWNA+T+Eg73ljgVkMrmzjZbExbjGn+mpVd0H79filO3n3mTdJ7TAK9A4Xvrh8K78aC48PF
zgnrvQ0JqnqfxztoiBjlCz5PHzaBVt8/VljC3MpWUjSEOsWx7ZjaVeoeuxLyrbsv85KMPI0LI573
kT52NCLDtmkRisyQOqVnhAVlF2NPn14GNnS54C0N3tEVImrdeNjLAdLggWGw3LE14MgbsfRxog/M
W96KE+6jQs+KteXcBDTeGQBHVyEYjuFfNW49/scellBxDJQJPJXXFDMEMa/qRsU8/J7xKNV6VoI+
4w9cMq4AukcP3jvMJWjc2UUzBcCXdURfOHvY+4swVPZ93yY3EYEQAeAdcG+Ke8ZdF939nQZGWtUK
khhMlh5ZdXzXbu0420ZesCLNKPBUaxnbOFSPUsDP7p1XIyDN93WxEjjl2rZuqwdSRHfutJabhWh5
DM2Q0877vzqQB5/ktGjIKf773lIbbVVbSMxLt4AVYTWrr3hh7XKvgEIB/lqEFyW6T1i+flghHH8p
WMhf5Me2SSGJ6mpbCoySXj0UBx7T5iP0Xe+Pl2DUvaSJzoTwSeC6nf1m430Ka5CRJ0BR07JnlIDK
CZSiBXOYd2eNn035P6HsvHZ7nM48JDuFErbDp8FfVLD/EcdR3D3faNT/AktT031k+YVA+OokkUIK
Bl4DYDA1ll5/5+nBOKTn+fGc3oCWaHz1HQE/1wv36N0RCNz9egPJsXhJT8CR88qeKL/KicyV2g78
EGJXipJSUMYtc44CeKE+iRpe7PIwrxqC8vL76NdlRnynbTUvTRZgNsv686nFDQm0m9mqBCgmLr2q
xHHvoaanZ5niZLktXSVg8c8TQ6oHJf/JQ3u1D6r5c5zOWotu0Gb4HLFIUSPLiYiZ3WBXuQZsWpya
qYY0iXcinvqGKWZERoR0BkL4rHiVyVwwsDYTX1RSgA34aevjrw82Z5NkjHl41nlcbL7kSx5E3jMq
g82CMHSzQkh6riDaEqgydQoLx6iXEkcm5IbyQf7nkzbh+5e78QNOq9oCjYO6M2nQvad3oufAb3rB
i67opzdFiM6Hat+1/K5x3jUH3zIax0HhJ1cfliqHd/IhrYXasZlAH6DHkt8HGrbg4SgwHskjnOwY
jCkB/7BZne5/Xwq43nvQoEhKVQW6+ct5pqKk4XFNi9MQ77317wMCvnPcHTEjpkcw83TMaeATC6Ss
obSiCpeF3H0DlrKM0jZNw8PcOLXZIqiArlx5AROvX53U76xq3JMq3j0s+IkX+CG6nNrPz3PODO17
2rYps2hImzM5Tqk98pKzULzTIOlSuRFuAvx6qMaC+Ii21ZmSrwvJOT/AL5eE5oTtm34VdpVWHu68
Fzmpa1oDpfDdH942sqqw0SQz6YhQJxa1K4g1yMLuaVZOF5vrQSFuoYp3/FeuaMgDj/2e5yg2FOiM
AHjbjqqya+rWHTsnasnjA8mz6TE6/lVxWfocMwZZjg/mNwr5QPF+zk7iVhvuZ1eUSLLoQCD4NBSH
NwRvVvPabk4N18uN8q1Zu5S/Nm6G97YgYUMmwvgjzH2tMb71K0En1+fWyASj4iujBWq9vJaBpNXg
0Qn+kczDtNZmoui2EeGmIlCmTMJITtsRw7y3rKkYE/tbkIehhWm8Xjm1X/bMZ+2dYrzsydtxsSt6
JNvYTqLqS1pzOAParAqx02m6o9xw19s70BgptbSYqtaJpWvXUIyo7jIhA4xkwHbz2XnWDX06ELgJ
jOhpKHdf0pg5jS7HQ8KRWEoWBjBlcQ8LUvPalNqIZy6Zh63GJYoUhFsuogURarN18K9HCIJ8f8eH
HnCgXeEvHl9L4CLhRl/oiz0MgeE//+r4ilwkbKzgWsl+lY+neht9jKimmT9e+XMcLVY7uv3e5X+E
4uNzC1EWS1pvT7Qn47DFxrqzUobv0rZ16HcT55G2KTSPqBvgGO4McuQ9BW9odLzQfyVUbhp/fW8u
hI0CK4Lb0gV9N5XS/tUuQQ6h0m+vVDdDVYpIvd7EAkPursRiUhj45+UwC+pyAfU5FI6jRSuTPGkZ
s7dxXmYEWKwzmiyQQbdgFjhHhEPxlYZ2NwlDtP1/KH2L84CNn4+4lcTCeaFe5fUAJ69xLRUZj0j+
0Flt/1fQmLY9HSr9LrWXjOqcsvtYooffhkpo14MeSek6W2kgMT9ZE61a6zKHQ0gipZTZND5Mv0C3
hAcRWHTtgQxDi3xyUA4R3AnZEe/S/a/1sNei3FksqF0vYZ+U/58bRc5giD4qyILB4nySRtzK8Zdm
0YUuqpDx75gD/iGJCCwL01fGAPnT9omnoomxPPgBkfYuAAoayV3TfT9jg8hEpTYm6X3XvRLfNV2D
4m2pDush2BUdkncYkPgthGSW+v/VDE5Q02//ecxtF+4DJRZVkhYnczJ+WOjq4wlZD+YzgKXKZdcK
S7iFVRwy+51eSbtXQOh4eSJfg0JN4fgg3KtHb4nmdylbuvbf1Doy282gyB+Q4Y7Pk0rR8nAlnfLg
lcQPtyWq7Cg48OKdvyWvkjxjN6MXfKVwOIcApZjkYLNsK8RAEsLznIPT6+FZ61rC0/F4mq3LL79M
FXh8fGrlnynCbbE/0zWiJEuxsFOsM86rbrE+yfma1V0yoFRqbP0z55ctJLtI2GRbxulAUaU09eFy
iaKy1kyBm6XXXDU1g1yktR8vWMJkYdSjWc7XY5F8A82/obEhWtC1fROrjMIqt+l0YeqQ4XiwJpFl
lk9Pcbl4q8oLW8SzBs/cceOPdvUuj/3JTW21O8Ianu9Cun+OC79i2pX1peWidI8Z475OjUu9MQk2
mLAn7oz1VEPCubVGXzhMLmtV0hGSJh50WwEYUeVozR6uUieOFpziV/uTKm+vUo8uqgno9qLkUEN4
Di8eQ5kdgmO6p1FjstkeT+DpwVgLq0kjdyYBXiY40aJOMkNFNoSZ0JAcotgdx3+Czf8YoR5ohgDq
fhmZuvJRoS6Aq8ezXCfkVS1Nrvg54rI63isJDJ2h9mhrHohVLJJdNiIg40EbfPh46TmRbzlqxBUU
lfcZocmLE6ZAN4HEVM64D2PXHA3rjfQqTL8ofgmmMUgoEIvJ0XesmWBjDXEC1Avx+mSk1zZAU/L5
s3IAkXK41FBrGNO4ltV8zo7MG2U/47i6LmYto7nzSsH5r9fHwfrdzhoWXDVNgMc8Yn97I7gYmzhz
u7GejiINZSnU/aN14TxwKEg+PA3/g6luzi3YtUuNeXg8JnDdt62UVdgPRTLQV4Bjm2X4L1hRGfTQ
jfVv/ZpMS/f02UE1e8pYcGuJU5aFeq8Qx8zHhGC0ncL6cMVpx0LgK/TyQMEU3w/iHkwB5qaE0OqR
cUb7/UNxCSEbJD3fJ7AWX3W5cURlox8uST6pHS57ngwpPWLvhgncpInEAlstQ3Uuw8MRlvsMaaHU
nv4eyQTQgQUwlptKwpWvvnZLABz8A/k0+G+GonG2XxYs4n49AanV/mSd25/ADXrrq+Twi+MYsIfQ
q7YWnekrtQujt2odFg3OUUzyxoHtd5xjTS05v9RmEijoPqbrN7l9fU99HitRFrzUVmRk+yYytxxh
7v54mJB952NcS3bCLoMOe4IJtB2pPXvFWukmP5quW8gB3EaUeIG1HMuoYb/yVztaifs0YViCSMai
zkV6zT9FdXuNkoCmn+BS3glZ4UteYAhiM563WXehWVWbELzE5eGxRKm44/vyxXnPrKW2xlX84puG
DnIYDS88sIoWMR/409VGpmJPL4DqWhajv9JiITc4yhVVEg5XPlBRgSSsvhj4RFLQzZ9eAn9XH3B3
k3C0/+RrOlZjEojqiAO+9voi26kUaTBUzmKr71DSS2a7JrTdvdg/hVKGfsBi2+ImqD7aocFQp9bS
+FK2hj2+CsFUSl/mFdRL4Cvl5Mx5JoGa4dEIRXNp4FgKx5RH9wQbmW5ZsWcKQ8TQ9h1RDiVqL4n+
TXamZb/8teCPUHi60tLU3FeamlkbSf6b5fFMvGdRbFFqUB2ABQk4qycaT/JeJ78nb39Sbg4M7H4x
WfVQjZFM+D/hRp87iMIiGzDXGbmW++SyQnXj24r3sh8BebEq/Ss7Uu4rgvjDhlBfycBZfdqcOzW3
rsXosFkHjRYnvECVCFF2aEweNm4v3Zv71+kiBHAIZ7J5A0iiGob0dVX0h7jC9TgK9bMi/tf6JKD3
TX1aug2SpAXHoAjT2zd1/00+qnZVjgFO7Ubj4bls142y0t/ZvkvLOhIkvz2H5YBdtAUPRH+Zbtz4
ApxNjqwj4Uuy0N3Y4zhqlSsVlhsrFBcm3c4B+Slo2wxEeIslh9qJ8SQ6be95MgZDi5WaorS9C39t
LMy8PkNtfKmT8B6aJmr2BjbFqArkjX3jDjY0GXZgsZOJcn/WsiY0eWHDOe4hF9OV2vaM1kmD75NQ
S6I+XQ1B5lkiVmsuxWrLfW1e+d1QGGwN3bDyVdke4XWfGAfI5wLKKcndKtkr+1KanXoRgo25/Blg
prcztwd+kuBHk/QDhSLGBSot2Czw11IPAVgayJSkVq8kt+ne6fgZ0+SO0jVSKSM/WK7LBrKAlN+9
ZgsqDE8wyAPO009kX4dHLJ77tmBLq28Fk4HfxJftVtzk+VQyp9R9fWwP5U1qS7K23kKaAvTBuWpP
gZxg0zwtAyY1douGk0NbIUQ7YD6JKkGPBFDpt2fB3yzknTziIMwKapM0I6h9UhajiqoIdJFGnjam
+2KBoepCuZn6tV1OhtAbXDEw10z4zAvqWin2AhV2EEmhkMWOcIxjdVeL1AhlkiMFoJ1kRuXPLnIl
AJjt1ugVEY2fTWVUlujLJgro9QA/mPqTOnlqsxJPZYDi0dWJtkgAKmAco22WZV4ItngP0C94jroM
cHMoXpWYplCyqVKpQh8BnPwjqzzjXui74sjoD6rqo2tdWvXwLdkQ4BttdsSNRn9K+pdLRB2B6g0r
234RAGD6zM6tBKwEEI+FR+aZk7zzjG0xJ4xxySQO4++UEKgwMa3dGLOiGwctEP8dpyD0jweDMuXq
vlxEvYlfvJiuiD1lQ2ZzCFOjjthpUiiZYSjJSyRrSa5muhaZvD1qqhvfROQEDqgkgKNPZPDWM0gp
zbku6pivXANCljpl09zG4cDTXghNvT/wjC5w0op3d4U3GO/GJa2Tw1XBwxIT7eeTlyvB8ny9FXOH
JIWyPhS9K9WUkYD4LAsutAzQbc2XHFlyOkyEXK9+UKcuoHrMSO25PoEIxOM7oohfbanR//uacF3n
h6OQQB86NqxBhjzv80AiaetrV82KaGgBkOOBwiMCiuTfMs6lZkCFEZqzRMU7jPhg6/RzJ8/WIQAb
iCvLvpjKlUrjzVyb4lNKndoz3F6FePnF4D35GSob21yyuX7Ac1oQZjffNJlk2xeH1fRFdsuL2lzf
Hhlw0aESH5gF822XSLSgBZeHy5BH9s8Ea2Bj1Bryq5o8VfnMPuGxCrTinOYGghS+DCG0XD8zpNH+
xNZfAWZgNPLS+C0XyVWzn2SKCW3Rc/GmylaoXJ0iSx+0cFWNvFVgP8QgWfcEg+O1Tkbyu9AJtgcg
auKINd3X6N4eeKWO0C8PMX0FQAIr0ZdZi+VYGBxQ+pK1spup6jHjo9Ry0y3ZWMNzg9CHBRsZvTmi
/+uGiRlfcIz0zN4uxZhkp2VPN99/BPPTmbf6rTkGes4P1dpL/ZQ0bfwgefl9/ev6i26hghp9S1oT
b2QbETjIYpmoq1O2BrN8bZmxi3vy3rR6/OWl4ASW2xNJCt31MaXMuNVaQgcCrMF8h54do1J3FS8u
NnVOZMAbBb17nDEM3dJ4LaUGvc1oZs3xZkWYJEtS/NmJfl5QmDjm2IQx1dNphJ8YubfE30WMOPDj
giiSlwH9u57vrJ7Cz+Fz3oAAywR+GYAl0fJOIeCa57bc90RAHzGudcD3ytxkOiwI2f9rb2O5nq8n
6JrtiqVTDyO2m8MB7Msv235C3uHtAmeoQg/fKGTVDKeYezb7Lk34vagSCBaH5k57gqpk2kM8MOHE
tSrcqETmEqTsCEmh8Jb5rfVHIwX0vfZjQvtWfOYk9i2qU3H+Y4CuHz5hCwElSYIOLHJYA/h2FPH+
0XFUCysUDe8pfMa3OcJVJ2mHZ+a6VKxLQqZZ526qkGa6GWijUjaMmI/cNtjoZ8QjUz6mb1zqHrys
tnhH5cdS9cRG8keJB7ZtYzw4nc4GRmbkx3/hPFlHpOqu1OfzmAjI2JoFTJDVSqnI4PF+mJ1XOrcT
yb7ZB40fll30UjA5O8W7wzyO/oHGCi9e1Ki7LEJVI8mCGNUQoO4lFWwCuEZqd3So27cHiMN7p3CE
fDJKr0nN+1jqemMcRAsx30Zv4IePhYK+GaZKdxAH+p+pM8qGA9MsaXPeOLTPVmFLi0S0VeFpk++a
QULlrxnYhD7pAPwPhpJ3DgJ44w8U74oIeFkTUiGAeFyrzwYsakkzoETBSiO/t6jRYeisTD5a7nlt
UHYbi/utat7KZ2Al6HvCVmnO95ycwZSwyWwbTUAynP479Mz/PI/rPgPovb8UwhPM8++MUN57pztW
5Wcs8wnUvrANot+1rKqUGqaUWYkMZFiokZLv55vqxzOushlc+IJToJ8f4v5ldLe+jAPc6SIKuwjc
kj8u6Q55ain+9bfx4saQcMjFBkhqdCD0oTCTeTvl2MGTLACl6OMnJ3PRLzbpV78JxOOP1C5VdhMf
1bz0PAV8esZqFOYEXkO2VZIS4gs1JhES47Nb8uUzTygMw+7oQ4TMWb/MxrfhDBgGV60AS0WSnX5F
neDLjY9mJxMH5CHmyJK8+IsL7EZyYOgO/rDIP2wNjEanlVqn6uoJBaF6bsYEDAkatmnfyE0CafU8
ngeTCWPncbBc+SiMH0Zi38pPESUfC+nkdAiCVG83eXtGFmttY4JrHz00Kuj1qhMT8vzNPH0vb3nW
xBkVEWHdAoAseiNIHb2g7Ll3kVgYh7ettkM6wPF5D8+D4JuXbYg4pi+mvs5TOUsKeCNNlQ13A1HT
ei9tM9Ofd521j8E1Ph+6ZmLN0naY/KNqgVusy0wA9zOxSADR9Ybrt4sh9wXQGSogMwE2AmyAunIz
pQLSUc8T74yMztgxZnt2Jl9GCmiCsEwwlFMAtlHk7IkcIl1rqqLlS8VW0C/n0AKy/dnkwkaTcAT/
yG/ybP6t/t79+bpBfxytzmkLKQ9cv3LFvb6zLhC5cmbPp/+7xE/9dIiJVIcs9qY5SM2+6kL/4foh
sStz2E1/sZ/H7YIFQ0XKNxsQufQCToLMzNeOeF/t28HGv9onddXDF9m+X7cmNIGQlTijDXYWOry3
PEF1waiWYhupLX5m0aGq+TEzA0l3y5WWrRCeiqZZx+Ewbm/Z4Ah+k0DkIy5qK7kNC4/YaRbMbp7C
DN3eUwyKW0XwyLmpV8LB6UjSrNnj2HMy0hcRqTk6XKxHMUN2KI8dJPuMJg8I88G/set7o+RjdQux
HF33f44hX2jVmU5z3XThuwANsy0UoXZrmJGfAjRLXhFjWj6dIKQzqL2STflhPA0MOzcQckuhRCvV
+PqV4IoXo92CV+rusqOuaRy6zTYloopiTYTTaO4wy39tLLmiuGF1E5MLQk9fZy5u+X8WLSl6q+yz
1WnRQIRg/S2iW5mymmK7Q1Miof1bPWbqH166B35mx8m6A8R18W56SZdsD+X/B+AYVi81mQYfY4os
+5N1CEL9e4nQGlmb3SNJHQg5zzJkEY4MOdisYbtTgKE4vw1FdQSRonATNbiPbQI7Kibvy8S0rxS3
nFq4I64r6bKpiJ8JSqmJYuLHZWFzGzCMJpp5TgVaf9dg6OqQQdNEimQ+wNDwm7f7N6NPj/YsgHq1
wvXERLSAR9zP9z6nO2nlgPwvfyfa9a1Qte+thDXAlxdb6lp2dKRC4BpQA9tJwvA4MPuhJLQNRkVo
WbkVF36FIBvBkEi+ZjPd0anANxp4nk/xOdAzaYLC8SDfY+fkTF7BGdRlekSxcU6332x8h2RPvxMR
qBhXkDt6P+POlxLTmNA44vqTjPxrNJ8I+bOkNclt4uUhnpWItlwBZfrZKr2h1vtr9ktfN61MKVqT
pmvuJMbqtY//TQEurTEyDob8X+u8mlS+iJ1t+PTXyNy8Wf7gOYLtDvWQBFILFCDZ/2NUy65jGjbi
DRBJ8RnlmMXupYvvqgvAxR4Ip1Y9KbQ3WUOwWSUyqGOW2xF288EQPJsMyQNxZLiebgL3Cvqf5mjY
qQe2iOu/Bz83YuqY9Gm/duRAi6+Xkmavoqtp4kQgWo2tz9jvk5f6/52B0yC59pm3xHt8D+T1Exjz
26I7stTEbYpMx3LwMvWazSBO/TCQoc82l8v+piscxg3qUJFR8h97wKxet/sol51AQUFTnfhEcnOY
cCXMH6JLxBQRgRLImsaiBIpKFtlEaimVos3PhTU4n0wecEihYWx93FcFhe4HCkpLOHW3L4tiTKnY
bR3hm8f2y2+fL4OCloyilGWxtioVassgruYxljjhp9Cn2d88CSk4GNnZo3oCMuvE6ThUgYDgPK1F
2erT0WhSjppy2Ki4A09iP/uVnriBkeFc+ipxih2KuICx6LW2PIaR2oGwfYPBt0jDyAdzx2OVf/QZ
BDm5x+ulPuIzFeu8H3FAcxZ5knT9xCXq3LNxkajGgkk6tAwlV5e+GcIk1Z5wzyjEITGGgqm4HJqy
hqg1G9m3MTzTVsl4wzkqHgdd//L0RymGIzbA56IhdVBEk1dafvRyB9ZlOX/Dkxa52CO4Jq5TiXZb
lIUwmWRHJHThXu/u93wdbAFFMRt2ggCh9u9sdCXXOaFVVbfvpamdXvKffauBLVY9WU1EziDSh24G
cms30IBnLC+7IUEyCE7Y3/bnLOeSO06+/7k1Y2XRkvdArNn893VSWfbll0zfkTD8GJi8gytDwj4V
ee1ikoru8sflSQkrJMubg2hz2NWQYFeVI5/+9qFh8cAhZj7vhGfGVDd5LUcbrNlHCoXTGzOuNWKK
HeePocxG5XLTesdG6ZRaRBVes6jukLYkUjnzrkUsYlrx2pqJTUE9heo/6VyGjal7qYw/vUnSpLZx
Uu4qn/mn1diZHrQrwRiKJL3MQN90y/45jHSqWgPJ26EfRKpQknlL+FqAAu30i9mHFjnig/VBU4rP
WfWyei5kXbmpCw1h8AVfTDi70RG8ygni1IEzZROSuT8cYB4bWI0xFUiOdOGp1aL9vHA2Xpla/nej
RX4GPsL9P2jYkf9wPPsGc/yhHfmmN/t0vLP3bvaTKderC7/fPh7cLLjcvJBBPFCWQy2AybZKmInj
XRxNEo86KgtIfjDv+fQzXQxGUK1ZfgWVrbWmTlMyHiTeVClHFV41Oe/C41s6AmMIG3F6JMNZ4EE/
E37HJEgyoOzZDqTDsDBGxPwvsVwSdsSi5FvviO2iJ6PgrL4W1vTJ5dXJqMUzBx0+OncTIieL1pZ7
ZvxMDbmV8OKnFpd8DH2ufbGkxZYs46SokiDFHLo1S4cJBsCV/pjiQtwlaJgfGSuXeNkckoE62u+5
vlsJPZRbVl+Y4I+KeS+aqVh0Z/ogVTvM3w0BjNq3jxkKOCVWsB/lyinAK7mWFeh2h8EH/01gRW/Y
LLwmMUtr5KCkgGYJ32o55IWKpnUiolU5FiBvqmbuQxo3jwq4LyLGTze3OzumtSBrIjmbGNOwLEax
1m75XuG1kHf/kx3bxE7NLNRfusJocFPgmgZQdI07Ngtfce+eqFqlXNm2VeP/SnBEp1bJDqsSTh8p
tkgFEY9o1pc9ive1joZYWydQ3VAPCaAt/kd7iBPVPqARny3d4Ya1nYnyRTVB9JMK/9vSQeYWqAtl
D70paWBgHb1D6fjJBiM+iJtiuvp6w9PRaDe+A9g6wxzVPlnCo4vJINxSzKiDBZje9jwNAPgUk/7C
EiLlK4oXCLh2NNQ2rSbXhgttrhl6kkG2NQXsgD5ISt51AYXU/xV7ZNDr+slk49KjQQbXSoaOlC7S
segeeyBqKW+LiaF5zLXX3LHc06kI9s5UJwCiaApqsPwXbaeoKLAtT2sBVSdv52ndu1Atzv9BeCYS
+LfitBtYC0a67pAeFTr+78dNs9XZcW//M4rEw8KRaJ757IpI6+lRLGrKmJ+54zsCCL0ZxKYm9SL2
btyvsqyxLcmBq+ee978chLPCXFKPpGh84HiY+/0y2kglvlbFjgOBGHUswjvRvYuWY7b7rK801KU8
8J7xjh0Hw7qFfdVhWBxspzWWFDhx1LgQVX60ppkwuU72PbyeVxCk93yE5NJo5FvGjRAfCug/QBdF
vdQeeck++4s/bjePLN8vfiX/7E9joG6FYPfJ5mgYk5uZrI99qCA4EvHbUL0qt8+7DCekkE2Sf4JE
FyNkvkM6U3b5lfE13jij0ws+HZGc+S3sBov58BoQ1HBn0czFoFjngTbNPN1474owsoVxRzgc5fDJ
xq4NtjjCJB66wcsYZcFhUaEeGTlRY1eBe0YGKghFhgYMjUPNfIQI1gqJUxNs9cmDWRGnSFglwU7I
HLlL6txoYeYWr7EfzwM1XklLXkeAb4Y9DfGXZhkaNHu94Vubw8oNsxBvmyzA7VEdeIWxCq7U7ezK
6So/xxZL+4ZZ7Z754NLIH+B9aqJ8E026NOBi01mX+eJuf/se5JeEESlTdYglq3odDytSsUolJhm9
Ymy4ACvAJj/IwiQnqYQm87V0B97c9vSfXx9e/bU04oJqIJtLVWCDacr7eDGd6LMM4s6X58F0AdyM
9HvqqHgclIZ/SJ+vot+zMYcSLv+FOu1h2sYAfH8nK46z7YJNwgazlRuWOAaMfVGxiAoRzzFZOavV
LTGgd6wel92AcnFq7Z0cIBrNMuZiCx3OqF/OwQ98osyImIJwBANHrWLveKwkXmYQy7RSoJjlEOR3
b1Wzn1pOdhqaWUsZdr4c3xG1BCTseARl5ExEjbics5PibvtDynjZcxDk8hRENgv/tpSHnNkxkI3u
2qF4k0B91MYi70+DuRKZGIz6t96TBjtD+zQI/9jA2RuO31HpHE4uVLQZUcGKlI5KK675ZEkVtw6/
kPnn59EFjZBPeosX96F4839Av+RQL/dZ24f2K6pXTEgn6b2xvdpYQLzTrFD1lBsx/TlYxvve5Bvb
Ghn9yrLbfq5rrgbj8O2m9HK8TGOfpotaqfy8zi9zFeKr3ilNNu8r9P/y4vTwQyuZJRhEenf3oii5
zupUdQg9tdP/kZXaNEaPE76H/kWmYEutxa4vDEawLr/NINfQ3Mn6ypXOshQVCQTqEkZs8wvgP6To
8ZpSiGzUMO2sBx85+M7O1I6jd1Fo0BYMjpe9ncQwb9wJroG8uh8jxwUw+WjWyxALhGGnyVbMLSV+
Z6NqSW+AXe0eJG2PZjnJjCfTWn9sR6IwDpatRVb1xSYJyJq54V6LKkyUWhDx8Pb6sfxs1h7wtw07
5j7CAtQ9Mxx5/27nfL//dnv6ZJDY5WBaWZPXU75r2wEOlsm2IBmZos2vu5SxPH+V4c2K3cKHvZwE
rQfqfHrv+XqZ1M5zlCULtskJMMNGEP0P3sWJSy0tGz7d97pVPK7FUH83dOvWLSTM4a3K8r42e/Kg
c/AE6FWISw/g8mNMx/3ZbBM9V11Ah+cgCl6OJx4641t/kqU4UW6MplcMNuyTmGGUH3XFv3RJKfm8
yUTIvPC8HOF84LANibDcFZhbTXirP9MeoqLMOu9nyI2t2L+/+iZisVYjlKcbI4Ru8TUqxYeMugQ2
IMFTvq/TfL9xSzRL13XuVR7YstVILAPN3XxetIBhOHmafQV0Szfcs+LNa4jRMkrSYbP+kJDA8VMp
xSfEHSCajd1US9KENR3mFgSXrizWthmHVPz1s3sbRss+pOs/JtIe8o6LTF96BplgDFSNd22sVvCV
XFhrDkVnXg0MuFtDyJ+KPqaKba1IefftAMKNq/uUt0LSTG0X8u0su9qC0hFYYTEnJ0ksJj3eI0qF
JtjRUdbvf1mgL6dmCdFbiFIE5nDUDS4gYUm81edIIyk2hgOLBPRCbv7paTVFYyKZzLWOas1Tnr9H
XHwPxq050DXIHKKiUBqA5hNWratrcPKint7EkelZy6nSLBUdXCBwUWC+rVdiPnzWVXGV0KBCt51k
1cAMeSkxpY1usZdqU/HDQ9uaB0Kw7cJ1z3SwNSDpJXuD+mIIpffv1W7Y5VJT1bj7Kgid6xPavt/J
/v6vlfOkXHiwcGN4jZHcieEr+bmc71AZLaX9fJaM96K980DzpU6uNnCocWpuz0z9qqy46fxGChzC
vJk9mAv9pGQQ0dxmyIkGGRpSMOfoDS7ZwSF5+WtWuyoEpF1iWGf0VWE/6i/X7IDeKmr7ZjbqQ2N6
cMO9PcL5+dIe6jC2DscxhJOv4jFBJBjWQqU6Tf9EXvSAzzs02hfuaLnPtg5/z5Oy0Mmu1Cxvs+4f
9vSDqYjp988ZZtAvr820pY8a2C0QyMQcLqbM60Jquo5whMXDT9DppEr4V9eOHoLUjz0vOlpdGXTU
j/RsKXxXjq5h1a9ZX9E3rqzG2+a21lQxa9ETgoBI+ckBZZCcfqv7RdM0KCnyfh3tD1KWK85eplb2
uYDkQ06hFGauNlK8hHqKFC8srWdD/NVVnSujPTcQedoThoo4hkD45MgmlkkjOob+NE4d/rBjLFdE
7rjrANWdsIKY+GM0drhsYpqsLwnM53yfjONJfBkTz9X+L3UxKbQ3rKAJjuviyYIsoGwZYDLysV8e
VjKNmaNHKZA8kIzBth3GawuMzEs/Keq1kdqUwJOgEanubSjy19REaBUMJN8SF2vPIewUArBf0CFZ
0pU9WFZOa5Qe4IECPWGuvkSGyapmSMf0f034DRaCWAz/RIfXNet235w9NeC6yQV4/Tird42IDfzu
J2rDasxIdeZ0gwNQzr5rE8XXBx8LZSL//cypODzJQESMOYZEO0pA1xv0At5ohl2iKAmUdW3IwSrO
M6VLOJTtx5k8jf1iZPWpmfqhm+uzffZEYQ9rKbb0Nktf+gBNg6CCSgss7t7KbfpfehqtdzKnDwjc
K7Bmr8EnmG8VJQ91ouTX2t5dKraLI62tvy7ce9T+79Ew2YHEccECBGLiOUVgPS/3j98Vo5z4nSKD
yzmqZcUKYdZ7cKeK+3/anAB5+t0ufTCOy7H93tKnNsNU35AkSYXb62wSZP7P1jEPz60oxGV8Sysa
ftIFAa0niRS5PMsOEDmX3jssoBCBTFEPM1UrvLv+kUG+IvVJ/MIt+MYKNCH9Stqy5nINczpewqws
Jtc40DBj86/AZKixBPlgWMtanjRRMABM4Z+W5NuWx1adKh5mgLnvZvv536a3itsCajjNKwEPMs12
rnucS4DEo++g+XioXY9Yol/PZW6JE+xPKtNRnBVY8UNUscOCUgthCx4i2sowazbor5mwyj7ZPviq
aXzi4MXf63WAozz0uHIMfZH0Pmew1gMdZWfyQ56nRVYNemzkbmw0O8x/kl1MMXt+M5ELknQ58bG+
P8Jlh4SbVMqT0m0fPgZKqlPEkmX+KP0BpNCMj+dfsZIndtHZDrstnxMJVuoQbDGwqrm0VYr7rF07
ikFMODqTm5HbDSSH/aeqToHVfVIb81CKJ+Tu5TYkdYewPi6xjgLRCmsRQH+dITQYwebjFUsbcnvo
JWVmq8/ZsMMZMkkFQBjMMltR80XMtoa+1hSqUjiUPThakHfmZnxrw2wr/3mNWdt5HFEG2EUxBLIj
jQJY6QF6Rfgx+HvYLOkKj9UErzaGh5C7bpkPbEnidIN/Vc+QtSWouhgWgOWY9V+/QNKRFFYgteEd
ZiQXhbiKEhFq6BDnQ0D9KnriSKdt3pks0g5rYDcLzyRB3BqJ2gBuJeSHTwmthvl9f+U1eB0ma13D
6fyTYo/+S3f260CmwsMVpR8EXNFnAVXF05F8KHN0B3V6UJ1Y5HsXoeovh9CrmrOOH5CHvW+dDsIA
9lV9FhXKePshu9WQIVfhFds3RK3hE2vY7uJ2CU5+X59Czz8ywWfpEHFIron0eJ4+chjGoYoBKHd2
F5/Jua6vOsy7yqo11HBBpiIiBqgUqzJkyDf1+WWtf824JlIMMiWDfQICVj+Gc8zS8OVkKP8r2Wzd
eCgkYyEagCGEUanye5JrapqITvEE2S09j94hQGmrzu3ZiykIwg1sohgCKGOtNnJKQMS6z6VxMsz5
2DsKgZVJo/GbrthZvR92iEfBGagUmBUBP5F2uTcD6zTje391ADIPeZMdbIUnoL2BM5F5emK9dCw7
E1OS2l8/X21GJ4gQg8ZaApkOyXtA0JLnrYEVF77s6BP0xdWFtyWHfXiWkCahWbl6A2S125JtRTY+
gIWmhdrdm3w/OIXg/RIDlTUQ2uTw2oPw9R+w/G1RLsW/2q1k2ADWHqDJnVZLPfwFZdfg6YnnpBQV
9ReIOLT2l1eYfp8Xuacemf3L6rKd2+4jF5xurTmvOm83VvmSDkY/37tdVCYImKueo/w96oL3LuZt
ToI9sXPRFg7Z5SOkLWOuF/yDt1o6lsqIbx88Nr9kHLNGMm2VJghGxeTRaqOu8NaB5kibQI6blwmI
PStLwAOPqmTXComQKAyoLqHD4JyV1+uNdYWm7jBCo2dKNWrJvvr4hjM6ZLFPP+Jm+diMO1noQHWI
oQSxJlIQw8mncm8SmTI55Hy87nF1E8HGZ6J8yQKYVUymxBuWjHL2Rmlvl/txsEd3jO7eL6sMWvvJ
rG7WhGAmFC3frJCFnI14nx4OXVsstPsF8PrwG61tGiljynN/AQKRAr9G4m+lHL4mgeFu8DGeVi22
aRmOtUfUXuoXDkCVvA2caEuq4p5fLAaiRPyw6dNvVCPKErwOGJYr+ei0bTw7gpRFxsfL40VoqRtR
zMJLGhOu4W39qlIDS2SJ92tP3pFLSKdLbAP4F0CP6+iJZkxRzveSVvlDjIJXABLRHjJLRlcmebjZ
506ESNlotx38E1jQBJOV1aeh3HfCRs1Ire1BPVjQaKi6bDlFSqGE/fEJVFj6BW7bpFDuunlSkiIt
HmCtylqu8TKf1wfs+8CI+LOk07AkCr8BbwDqDUGMrrJ3+WcGYlLBj9JN14ffnTBNI2yx7CTjeBMI
KF5bGI9UKB90tdKgzSkf9O+rieLoHqPGRpjwqBALOaZylP8j4Lc5ycfMMgpT/6cccNQg23kqgUnB
dt4JmfG8wZ7WLWGyT8JHC04lZAIkeHG0e49+Bss6bBkBYqatG53KvJXavSBPgRyygHn+9JW2p7Rv
cwWRTRtX3kPT5DZVLqiaber+5Fh+P8ZXC1lUzlgTrFlnVuCxEEQYorvJsseEEYIQ5dfMqbofZj8d
hgXSnODsAQIRQ1HXblgBkcUyBDluC03dOt1Li7SXxgb67tmetdTg4rZprTZ6eFrxanLfX4rLSb5b
BGat86h1qo80gPen42DuFtOwhbSPEP3d9Dl7ilycrGQ+hRoJL61jBSemfuUv1nxGOl5E3PXBunHL
Lwua99GBF+fhGKt/jGmogadwJSssSGmRTDncU6GDiyFu2A9/9FzIHWZ4fu8kgvfoZnROUXtFQwgR
pYA3M00s4h9lwrnBrZyoZTd6T5376v8hPlhRfWnuwSClRARAwoeOIWzXkO4mI7X4IOPsF1klan4L
SrtPmoxSAB0klhVDKdejtS3sO6YxHBEaJXK778LZus19kDt4+sQiircHs9s72bSaRajwd4xDCHwR
y33KTiVmlut0Z7pD1+68s5/roBgsfpG1BxgS/IF1vN5shlzWimHqWGdKXk3fR82mgQL7AcBWUOoZ
lE8pvYyt3Pb6ihBSd62htHljbZuK3vbrU7w0zdr0tEKsTKULmNvUDtPvMnDLJX8+t3aa9buDIh6F
tEvzJ9kJyLb/m7UID1ep7TaqWW13MCSE1t5q9U8hAYqbbK9UUgFXcc2P3e9bde0G6ELedJ36SKea
VosTKqsd/dtx4eaSVbA5RMFAPzX8rr/h/2VkWjddAIZX7WoDkMqRdO57Jgz75cK+44A0g3xaornS
wXeyOl7ihDaOFGS2zrjx90Dq5u60LlMr5aRPhg4dBm+VVRkYPAHcGO8uyI3375IZFhLNAICUWJIK
wHkQWB6FHSh7yjKaQNmChCXqaNtkLjl/5PCbK7RWJfQUIJSF/oad6rwSq/QG3Zj5qb9raNf+NdSR
fq1kmK+yr6oj6T5VyAysIzVCOpfRwtICQYH6TALAYKvmETP/F6PkruafLma6yPrBDnizgvkl8dXQ
Nhcqpa1EJqNvNKNeuw7yxr7e0xovVooxXsXIvLaF8cREGKkN0I60fLdu9sc3EYax/Vq6NcgKNIwz
+FsqX2/eZBmC4SX/ge3Ix47JIqGW6pVBI1Ve1r9mNbP1c111P2g8dlkF7JFgWL/pDN76yvrVFyWY
AGzkHra3GKsDNwS9+rUdUfQNNwi1JJkMrW9VkTS+Wq/Ll6Pln9oL8PwzbOmVTQ/qU3CSDU+gD6jR
I17O0uRfSDihCXlMXEw6LTFB5Bd1yDFX9FI5ZT2a9HPzzAj879Xh/Zd9vlDwQey2pgR0MC6U3m5N
YPI9umqFMtgPOu9W6x+lkXcYbxNMUNtNv14HXI0MvRuu3uLl2yuByauuK+tsw6fEdX/5sNv2yFf7
5037fpLd1BuJXhFUPVkY5XjPV/9gnIwk1cQfmVkilwQg0KMjmh75m7HVdH/8Ffsmup2/GI0jSvyx
awQEpol87lyF5E5+iOckeKHMIVHitBI90vgBGka2SUYWzUaQX2nBOmxnLQmHktz+pF1N5u4KpsWX
e4vE2ISPluK8Pwa7erEhuvNbbXNVJl1t160RRVjfuZTsRn3jc/umUzuY8uUcFWuJ+SWEev/CXX+o
e2X2EZhMgslNg53jQOOc3kI1PaLvk7WDJqzk9VMgQKwVutqfHA837Q9d6T0fOJPetPIYJe3Ko57c
BKRqWQmR3c7d220WmqjaBhUZ55Y3oNUCcxZHtQL1IXHO0vcNsAkw4SGmHGSvkTu4faxAp6WlUSic
vseeORZ1ivWgNFOdfsuI26HfhUxs/Zx8iLmNXfOQ7C44hy5Jqo2SdhIIXoxHcGeN8222eMdg2AhD
az4CNfZTCbi112V3mUVJdNdRI8v9Scg8YfCtq88luAknSb2LIES5LnlyJJbZ+k8Wdi0jVu0LiEBZ
+ubJ2x+GVb3kf57tVPOqTn5uGwF/J3AH0TMX4a17kjuUECjMt5Visheu6oYQG45WKL+t/zoZdmSA
fs/nNwlocnYjrCOTsflhwMDR5D4aeF6zGdutc1FzCU0DHIkShYhKrcwh3X7ULeY/oIw72VWYRXAW
Mrau42ckyDaoh9JZSqC3tUAf3NP15Ya3wTghQ1iTrIjdTOkLH7Ye36xNTdR6YZQ4i+pRLXWOFVZv
po8GV+auLx2yyJBW+FWeiS2GxKSwmdefKFpvrqyjRNySLx6D1Z055VZnGIpAxIewQDKUT9hGeW9L
8Oqsb1UnRDkSi+5YFHRaRbnkRg7Asn8P7/RIs6RU5WF9zGgQpt13lXwdAvjZ1K0qRhQWWdNHCE9s
wnrXPc+zR6ko32uyQQrVJjACNoP+3IlSYA/EbCWdmoNF2fb0j+K5E0GB3I+bMHnAn5hhcFauw0eg
4Wm6Jukxh7SSCNaH+jubVCibBe+yJzmtxupryEr6j+UdJ4ENDhMrilmJ2+3V4q7/YsB84Nm/cci3
rKPgn6h8VdfZwFrpdB9ucCGNC6pVGFPadNxzOyTaqHctvVCHwoFoEtN4shnBOVhrC8IijR0AzjYW
JIdUmRMlW/58F/btBsH5L/z9XMtjKeR10Q/EWgZL1zWEh8CPk014M268bPNRka6WIKtcsHXGRYYH
JXf7IVtfCfW5t7vJN9F7aSwpXWGYlg1KG8yRbdISLl25TJMxoORqJk/4zv68h4HVynmydw34hxNN
xSb16ochHF84safMCb/PM5Uaff0M2iiQkh7TKSGDr+knrYm7sX6RUedoICuWu1uLv+WKr3qOjQAW
y5tbLyCWORRGhv52TjYGJ85M6yn2J4xcJMwnh8L7g9Gc1FMTvaNUMcdOnQ8Rcsb1xwuoKEgj8dpG
Q0PruDgRcZPZviPRrocb4V2UBP017+5SA3j83zCPC/zvd6fET9GH5vrvnb2azfBXNQSbwEgsw0/1
4sXRgjzZyKYyY/fR1gSyo1yubij4A0cP8bbM4IsiX0v7jNsoCwi/I5WStNgyFi89s24RxYEj/PNB
eSai8Gw3II3pe752gJkYb2kqcPaiPB5cDWo4v6zg2H8YKjuLG47D1rBQD0IE9/hfY+uj/+mu/10R
Nhw68/EBo5KcLmaAJptVjhhxobevbMCoeOXV6k/EKtzjBqwykoTJS/4jDiaMqnXvAXOGkjxXfFzB
FWWjVv1+S4hr7KLbz775mXIga3mOe8HarqLhvBOV10e3nwfxsMXxshMaGF2pJrRIp+Dzzg+U69G0
Kl4tmwWpwYuQaZ0H5WwXQGmDnrgN/UgTuDDTTbkriDOBfDxG5k6rch6RFgEqemNF8p6bCrlUm4WG
cRoOyQq6BzISj1NIgF6bkyUTObqc8+OWqeVZ3YyXXTDo0vYxkLyYWjL2u+XNaWJTikZ7ZoAKByYP
mkCGvQPOdXs3UnscuqALT7soYGOiAxnkXXYRVAqdLzdU4OACkQBTQCbgSCjNAP92KdxLauGM8gk5
0z1SEJgvGJo4S1R+Td5g1b272qKSYB6DeqaAoG+hmp15Nq3nKl+9fv9wtxnxDXo0SfEXYM/XMT5R
l1qPG0WYXGemVZKXc12iPBlgIuYiXCKf5tlrQC4XS1/QgxTbVBcjpJhOMusWGzWqUX3fKfuBM1hE
wvvAf7cID49Bch1dcF8DjGTBSKaBHyotL03rgh2aR80T5pQAfHcKmG2H2jBTXRqPDjTCxkh9pWyN
z8Viej0UzODHven8H8puVwli0olzKxnBnM8bOqvbJmR3eFhGRyEmgQ9xxhy/BhiyXSwksmgJ54uF
K50ONYYJGQOkVWqTT7nnVdp2GcWE/rghwtTxIhyKOY89zwOOOiJELx49N25z2t3YvMk2jtd5CVTO
Zod9cBL/lP1HajUBmgE2QIGszWWPjyH/Ixm9+fVGfyqX62KHE8x8Auwd5lw0ZW0WMjca+h3EML0/
6Z60OFVhKlGXT6soLbvErEhFEuxX/ByXtFfyf2JUnPLdaE3URsZ2TrZ81KNCkF0ymMI3OuHRXC41
59ofv/PYrwNQEDxN8QkaBYZSuKMTb8ddfI5HMaNPO2qVRkvWgmGUJsI6eY/NUf2uUXT4X0Y3cQ3r
LtAiTiKqJD21GgCjhBMsVthgBqmBZPO4bo05ceT2WIy4LwXJ85bUK9lOsHxhaGUOXhYT9RHoJkFX
08ex2oLU2lfhLAch2NeskilC+/zyAel/17HC4ewF7AANf/cAoD5E+hhrNFRHcrp8MMQzQqz7kpq1
d3kcLCf9m7yHrGrGBt/zkv0iCD7i9ZvNK8erbGqG1zvLpFywYf3ngR5phfn7RRQHeMff6VI4UKom
+mzj36blG7g0ZY34QpG2DAw7VYbqUQj2Jmo9WXw96SI46k5VbhZyfn33iCV4soZzcW3PZxaqY4bm
3+lGz3ZYWbGWjJ/YHNl9Ut8PXFPWZYSLb4tJPDGDzyJTv9bOpS/7yLfOh+TVqSSzcwNQ8iUtpZg9
KuIM6j08PaKdioSir6HLQYZ8U3R76yLpwGHY5piX9Qhehl37v6yzSL0WO7ctFuoXmPIPosuwleXY
xvDERFz/OpkyS4odZFEkIrR6z5TVtLCn7CTn+LTEXM/F+KMIHYGOQHfMqrTXIPNY/dNaFf6/Y9Q4
2BpmjIKCjbrYeBsJExLrRL8s6Odf/phtzX8/Ym5g/Rg+0JXPw2relOVPoUvUVsmCto8PqnAcZnxI
4p7HdwGvv6XDQw1gdkd/pakBid5qVx0phh/kpoZ4ZNjm2+OuMUDQW0UXSt/XLb2NSGMtvwKipNqO
Ot+a+frkvIkglSb4dhVuZ0fmu8nNgim84Ef0e2wytOG3p5y+Q1K0GOXmjRWmq1GuGgWoRgGMXUXC
n0VYGwQlPvaBBSI7y8lHTuevV2dbOWEVCj4cDsVW+nJFeFk/mIyaO29Dai9T7D8SHcmgEOTP2Q/w
3oz1O3rqeO5ClZwPzeScdjsMbrysGW50knFiQ8yYHS1mJHVqw5KQU9y0LSXIEQaxcLTRL0p8BlHM
k7AZ6HuuAQ6R0kP8QYeBqJHEaPKFN5xuweQFfPEOISbsh4i17hAGhgI9fdP6HN7wdGmFfQ323B80
fHW2Jima/9cWy2lAjW8m1UGpArqOig3bQ0WkYVcPRoSFVMBcqiudI/6OBmt1GXGofx6SrlPpAM8b
lleNTls+A4I9EviLN6/kmuDVedxyuy1Cbc19zZFRvTwiIlMezFEDbo7bR0I+TVSdOLJ8BKvop4qi
Bce8W6GuI/8mapYlZo1rpr3jWD36SsPD1HJl21y+dr535Q8JRXsX81xy6O0ZusNKdhMk8Dv3XEpe
lJgRhKpVbuZ4JyOTJhZ8pDawsUndI5SG5eEHO7trOcQYWWQxDSOo618uNh6m1U//SE28BSAipEqo
OSz2csJ2GFCjhPaEoHW0J56IEdDes/71Ys5Wv+Mm6EvHF2lIe4lt+OJf1sgq3/GyLNL9H8QSBygE
ZmO+/cNX4ABchdzPsQtfzdp94NnYGnkstecXh2Jmnu6upwd/br5ryl6lTHhNS24ycVPiHf4RVzX1
6aitTsLHjrjX4xLFmcgbCBFjqY558Xl5PKo6Ll9u9FhqXdQhNKH/Dx+WZQKhmk31EIbeIKrpOd3s
sAdMdi0jFtmqmTXPVDCiedJALfghs8Hq30Zop01B1GrBt0hbjTNhVtcydMTWPd8YqDzpCnxv+B9w
ELcQ8F6iDsR4o7nFn+JGCsJBTSu4YHSNAN040T0dErFhFJ0qn65GmRh1I+SW9nzgV1UYKH20yTiq
pZMg4JycFDeeMooK5OW9TNiNLC+3dj8l+tJFiqNjvHIhW+AYE1VwmPQlSgLxpRtTiOCRYy+dkfPE
newlE7O2KH7C5N4cddsZoHYqAtgBjShT2EUHVQJfTIcf98KC5mA4hdE4jJuH/u9Mt3UUV5UYAKlB
LsmKdfbTaDL+l70X+mBMkU1t/AhBFXx5tTy6qgz0NDRqshqrPRyJ43W6FO5G5bzWcdiwGCq+xFYN
wrP/X2DJ4uENC5m/tBPkkuLsLm11Ge5dfl5n2m+F32kbZtOzyQ5yVDZl+aBQgOc21MFYq2zZPpNr
UfXJ0W8YN/BYvP8cypI/9itFhd9Im2Hh71MhbwatNYq45lggkch3epI2phVKRIs51/BoptcAg5Is
W7uDGKLfZrYUrVVJz87TDh2OentiBOAvMYxGj9ISToQxwmftaZEWJKCpm1ft4o+lTsPBfxkRuoQa
sdYdFrk++7Y6a7C/HxwUnfGJCR6Dec4fYmRLB1GR3YhPNzsyskpyqu5jny4NoqJuxUVp0wlJswxz
pKh3GkTCcIttLLCy8Voc4pKf4lJQdcjSE1ybSmuJ8fX2dLJos2W/z1rzNMGogTZiLzpgAF+m3mIl
XawleDG7vvPpBYMTtF8mmw6W8ePpHLZ3dZw4OXbszM1NKh9Yn4qnGM3CSZxAb3EgrVpXR9tvUqLf
mi1D+LCFnhW5msd4PorN2CCnc592k9b75GAtfl2lO/4ZlO7VSg3lzBs0xzO+xvFyQpZ3vHMkV4OK
fROzol08SRWP8yllju/FnAM2GGdA4Mykha4TMJQOERwFTUX6Hb2nfbBJcFlxGMiD7X7SGZrRIw35
BORPs4GZza4DUT20yx+uJ3ZFuRmpTql3Ow755MDxmkkqGq1E6OxmwGebOQ9v9WZLqnPibbrEJuU9
OfRLHmFcSBi56gbDYWDceiZJEh8OhWPXd4EKwQkfUQ10ipGgLJjQw/coRb/Y6LPCLACsJlPw8mrN
aG5ZqJVOnJBdyYhN6RUhBnw/LuCvg92ULeYlDTzfTikeJNjH+kdyy4hrWsJHyv/qsW4KAdsgc0we
x7wdEL75QIuGv9CThAeFZ20cUp9MX5fH98ctY0T0JFE4CRrwx05U33kH4rFmdVu4KEifGh/v4Nb+
M3MZAm+Qwc1UFDRERAQzHvnmezoZmb/2TEakuQZ4w60WoHuDl2SikHrOSnqEeg/uoFWJX//eh7au
lAzD3uy1atxfDFenMzz73Ds3o9mEpI/HV3xo8OeWwgfgXhG07ygapzA7tcIykSb548ddTtAe36XE
ujpMfCbEDUrZs8gOhysNx9dlUpNsps6oMaJ4v4f5WIP6ycpcuWTpEiQRf4gSCToC7VQzKU9ztXEz
27zcu4qWbL1yKLQEDfItlgrEaUWmgQGvpkCHEnNxEsvxqrAYkASNiXm95/zhbimw3UrAUcOfVX9M
fAQ7VC2hNL9f7j/PctH3H3pXBVvzicX3OcsBVyAo4nfOJkUgXHhB3NsbrWIaMw0A35/GRvt63Bd7
Rm8R5Tq+VrpXSGtWXFT4sJV2diAL8Vx3gIG5qU5zzKym/AGJsfTitWSGRLYyHHgeOB/Ap7yXheGS
yreEqDSt/Cjmm/cj6APsWeIOz4orQbdWAff5JPqDOmNiyRzv9wbruX6OgAyTLva7eZFtgILuLrI+
m5EJU5bXXUwdApt/45hJWOl1JuXhOQxm2CIhY87AZWEpE+j97QjqUh7EcZQsoBbSppa8p3J0YQw0
RRhJ4PvY/1R3hMIclhJzNQ2HR6576lBrDl7yvWES4yJwr5TGtEybTLfPZR29lmRjUnZcCYVhmTPo
bEHexlVGvv/NRMCbpnev49mpYS9bUKqbzS6CLgPhc/fziTQDmGCluZpdluKMBSXcQR1LfMf+ivvY
QCs4JdNZxkOPliIaVGmi8WKUllDX0AyTcWxFlqvbpCmytvmEsY2gP5wfLM4ilRg1LoGWvm5D3uO8
ezuDjvOVTEgifsjjHRbJiHu3tYeUhc2vEldjwg/XXFPRvUcl9Vf2Q0WRyRg5T6r3/9K9J1S1E7OQ
MLh2XX+01xVmMmcQH+i/0za+AN00O+FaCid725Qp9JzJ4lVvBXc6PkRI6O8AbLJUaNiSVMVVdxuT
SF6ZVN8BVPyI6gHdhrykVYp22zncR3IS6JcS7f/DutWZdAMGqBVxXavJ8Qi5LoQ9InIUE0NrIvWY
AcMfHN0x3VfbK6UzBVC/v0+EeOvHwqvPA15udGaSf8jShzwqNPw8VKLk3PUca3Ljj7EOiFe6eUxt
RYk2DmkbMeAQl/qQH1Xo/s3FQWZ3TiUi6KA3q2nElqu4I1mpnw7Vxj3npkW1+JVT9tzDldbjLy5F
b0uOKCeNBGJ8BIWAg3lmLpX0RYo7d4J5A/jsMWtZDHrlWhugN0rRaW/t5cEpriUq1RXN/Tyk2MLm
GMnjFewLR4obaAzFv15ShLgsB9klBGoatWry0/XveajGoEErYAxqT+yQS2HMVRkL9OPNxKewlDNw
zgdU6evy+3HY0s1Qc+R5kDRPA+tIXyHo7B2cWhl5EPanIXQW8LnOcy3alFR+jDwnechncUWJOe/H
OZMSSlpws/Y/l2e/GAQNAFZheYf6Q8kUkSncKwqMKeJNAD1iljJv/58BsOsMPI/yeUfLVmJfXLOf
MzWtfOaYU6LAz0SxInsNShIh8pCDJcSiVeDhJvHVLoPU7PjuIiLbXD8vUGfRjLF6wulfgTFpyYCa
O/J/WB9rPOfvq5Xa/sk2AYYc81fiGlNpvOQEazda2Ut39+iHT1tH9324TUGMUxCabH+yJrFVVDY1
oLPpcVPwmbGPhiaJuGoFXy67aweJAqHKj5mojovVDFsIIFjlGaeE2jaVJpT6COn3pdgBdQsg6bN9
Twj+we5tzdtkUpITDfGsrFHoY3WOIMh/0mUxS9/95kVSD4Tghf+hThlNHoNE4wlaw/yLqCWAVonr
YEnzN+2BlkDveEoISXvmouVKHwt4PK2H9Xdj2kumlrd5HZLJYes1ZvmKQwn5lKPP2ZTGgo8E7Ke0
wI3ra2eKpXBFbE7pZ7mGTXVJ0FdKl2XL7di+rXWQXKiAQlcpY1YGjwEiBEYq5iJA4nnz08QNoaNk
bKJPfJge149U0Yf4D1ks/B/FigISApA5ZINU2jDVQULTG8CCm8HQCA4M8Mm2Nhx7aABeNKGMYhuG
GCZv+TkppEK2M+kGn7b+EQ5W4ZNXbp8o/gJMhZKZoSYHmgxZiKxniDv9ccxs0cugHT2/fPjtu0X6
gbZGCd7arUM6jEod4RupwoDmxWQyFUmdB/ZUtXDloAxiAYna2jV1+ZzuQ0L9hQZlYZc0sCttcF3k
bHV69XYatBB37SGM0iquGxFwiY5baTQuYXdM150B1Q3msrj8MVmjPiWxix0zR70u6aZFwRmq2LVr
B09RbniKoQInBrNjVVmZyA3+M6msZGbALhcrnya3i1WiyBD15F1Sy/SOROR55ZsyN384yCoSLA9D
H/h9nYi87x9/+SvB+VUcFRdPwxF3rWel9ga6b9+TOiIs/QkqyP6aYZAQs2X2pIYoO3hEkQwriJyI
IQZ87SBEVfFVNjqXcvL8seVKEgxgcCJTIcqN5Gb0IWsitYiSJVuy47i+ETppt3Meac4UQKVWZuQl
RY4nvWDA23g7XgH41ywYGOl9H/tvHQvdxczGn2Oo3MshAo8IZjAUnvSUqpcw6+s3P4wAqvM6TJIk
8UzdfnY43/aiRBLHoXWWVEOuSBYH8Pgd8U5GsyzWgNqJxZiCA8eljoESgyQxRtUl3atlDWbqyL32
cqOKHllsz7LFxs8pgVDuOg11GU/xFkoN5OnB+LBVp7JikO/+cgPPq8DMEuYePZfYlP4uOXl4lt5N
LhiFnDX9jGp6F8CgQSQoaev+ol1gQpQOn+NqdgiSqOENB1R8DqUfAXOUtvMGO6qqm/XriUmsDLYa
y0eRKIWEZkEYg//b3tKKXJP3rr1mdxpZ7/+fqDdoRHL2oZga5n2nLEY0LUl5I32Slg8XdAwkxg5b
YQGhf/hzcVlit/wdMR/GR9BfQoqNGmUkTMvR1u91EJdbDhJk7nvWAivG4bthcLXspvwJV7MISBme
L/7mymGtjCkwf/GruVIPcaALfghAi9qPysajue416M2/2abo5MtW+R5/KjQS0oHexCt762RHh6WN
itsYdjndWD4oQXER3N7qM++u3EG3BNtsKMQe3CHBQpTP6aKBTGT+v3JDATT1dYg2bk5jc+O/67qt
4ZGtrd5Ks/7dZbTJC6mrO+5HSuFBiVx2lsSfmpQ11ACfOtGX2HksRXHSnfwL+4yU+PYp9lAz9LNZ
Zt5mjQ28LIIDpVLiPjBNtD9j8T9l5topeyxYrndda28Zrikn+YmBCQs2ZpZl4XkInbXfcVWHMlWX
PBuRMdM2ecmdhlJzO12zOf1HaqERY3IRu4ppZTEaUghI5Pk0K7xOavGUo/VFuzi9PljtoAWSnnej
6RpYaCJoVL0Qm5vYoMd5Z8LOwentC1u/kqVaoHFs3L090hpOqWobNFXlVUa2UvtGjjtTj85AKHjd
P8SMiDwpDW0V9CISH2AXZL4ALzg4TDMSPmdemvMR+uQl82t9+1dUlmGpu2T2Z9HnvGbrmpks/m2J
5K4paGXxv16s5/0tMk4Wk8RWBn0x5ieFFvwzk+pOpofxCe5U2W33X6Ew/PJlAU9AIcnmzYJQs36X
Psl1t8P5AJ6aO4cOj8eY4JekSQh5kYWXAjgbuChRx82glbiKHjJtmn0QJboOX1jprZtdW5p3OLFL
oZZtVXLR1BE6ag4Czs7/FhenSjgahN67OfdSkvp25ordYqnr8H4/Ky8Pml9S3Ad9WrsdM065eD3r
AzELRDRV4A0YwBF2OZuZtVc2y9c4ntemA7uqi6Vwhc0pix82h51LKetlDpPPHPg4zpRRm/wuz9Hz
gCCauhyt/ZXaxXhlqPbVs6ufyKBuhiJOTYo2BRTKiS5bX475Lac6UF8QQto9QNeRpQPs+tL0pBqK
w+mWS6qupepXj1S3RitHvg7HS72/e4iw0MZqj2/UWKWjqCBxvZ5oxmP9nDkmbD5Pr0OjdETdzHX6
rsspKL481aP+VkOgnM9XZBB4s0fdX0ZYm9BME+366WSwJ/QBdE5Z4XQICuHKLAvWWvpzUNIDLdcs
EzhR1SP2sFmvljdhoXEbdDogQrCr9UcgPrCbNQSI7JL18FhyBoUpxsOqa0rpXwjKHVSCeVvKZ1BM
jU7q/N45qrX8m8Ql+o27ZRfH1xH0fznIZReh1aLUiZM6lzmVzVWA5s19wxuhnLoa8ZJskc7XDU4w
JRhHhZG3/cNREe54ChXR6OkO66u8KWwk63AHrdtAy28F4rZMzFG52v/bQYWOEZBi8hB/r6K1/BtF
dt+lCu4+PGfWFue5VAZb5cG8/HHZJ+QksjYTjSkre4vpDgiZLFiBYXmw0N6qqhSz0Q9d8s5N9DbK
iUjzUXVDBbQYYr5dKEqss2sMFUMCAC22w+pXWcZdmN6BgMuljjIMyT1JroD5Wak7CFcDlRDByu7B
iDPLA7rlvBFx2aXpjqWmUBDZIJ8mpILW+PT1vjIIx0sqRxIY0J6pBeqXDyNl23u3tVWFdKq2xs5n
t6981Mq58YECBqf2mBvk3JnrDJCDF4RWQwsJ4axpu8+66DL21WJEqcjUha2dueYpL3RTt1l4DV+C
2ugiWhsfAfrT/QNPk9g5uQR0FwlIVK3ja/qDLwv8ByxwGctLLW7VVTeS2pk++eniIFsARAPDMcUN
g69peYKUBacqDWkp/gC2mc14FfMugyOQQDE366O44wuH0DdGvUSH5fUbIEldY5MN52kWpt9OxuQr
7TIip0FqxjIjPi8VqPmF0Fyqt/tJ4PR6I1bGvb+otKDQXZt3Eeb6op6A5Lld5Tt+jn3EAHKhWYpj
ND/IQ+YBk1SsbsT3lDMiO6JSxVLHGYXEyGQaUdw7iPd2y2nj4netOn3vjxkefP9DOwTOA69dub7A
lmLNsd+M/OBCIbjyarRYjmPgWsLrZEJ1jc9RaYV7s5MqqAStAcAd0Y3fD4SYWSZl2cBZsUnfnJv3
YGSgx8IpgI4psYc45PS0GXYKyu48xSFIxgJs3SfHkEuAktFyceBDOJmVz6KWb8fGCxG1Xha0u2Oe
OucQQF4QJ8ZO7wqnrdSsvKAfseMIqIqC+ygTWsYKf6fFOf4s0e4TUS8baFZgUnSv/S9o9EVVx8VE
iDLepOKx9nUd/1TWhbwlZogI3M3hZ9Z6fB2UYpwycUNkpJ87lS4QL5PtCm/oWOYzUeHqygIK9hlB
3NGbiGXXOjFrxug2+PPjVLbsZXeq0ZHRbR5ehMKzELGnMVg2iojz5vEWlH5Ove9gctk2wOexbYhJ
znJO5cWNY2uVRN8nS2QTEcuuiIRL3S7f4q3skvUDBZthz1QDHzScwC36kH/U/5x9nQrFjVXtdNp+
mSE/tHJM/6HMO7s2Ez4XvNvLS+OCgyAiabB1vOr0VgjS9XJdbcm7KYkvqdOLMKLxcym2ASS5ZARE
D7vHjhqnuuLhNpxp3E9CocW93wMBXyUPRjL9KXvcq2d9fT8PawVcZMIRKQEcj4mz9CK7wFUBE/oX
1vfknG0v29eHFNjhv1N5v9d52PaGCpzOHGMjPniSJ705cimSwLZqXxHy91vmVkrDkt502fCzjdh5
AeOV7/QAKeggjTG7Z4B//OBkFPFrN/NtaFTD8QUiQ812K78EpY06Znw9ZEGqHmRv+1gbz343IITe
ocPcBrRe7ZnqUpv95waIBKcGpMgGhdfpNQgvdYl/J8GS/MBxHQsRbTYfVH29mHoR/0JUD1N4PweJ
0FEz5N99R/qLha4qZGFe0xPwGzF5RKMSpjM/sOdka8iYgdvt011cReS+yyHfwr9irFI0hi0hiJcu
bgGwkUBGCPDi6XjgG+JhkJd+wyJVOwLt7T0w6ak3wfsw6mRfcPazLsPy6GphqkPKJKwcJT+AO/Gl
pp8M+YgPXJq9Z+07fHXtEGegbgB1ZmJwX6hl8FGlmJUrmPL3hn8l+35HLKXn7XR06ZA8+9K18kZm
8VMc1VpTUZJrujLedlcjaJkns6fL1rOtwjsmM45gca/7W+Tkw5gye/EZKJeQsKLA9dIlq2hPPwiS
iaZ7Oi6noyTJrPae3gurZZNp1+FC3kwMU3EouiPplRkxoF/DArV5skuhtgx2xbJRS3j4oScPvuK+
y48tlEv5lfGqc2fXy0Mx/1X7yaRI2Gub7FMJcV/7xbEUFeth0vn8okuJfYsPC+8KVqd9zseMGIBV
sphK3EkADfdmss6jSR0qO/AbVeweB/v7p5sdrQ9CzADQR+E+OnHg6+Y4x4huPra/UqKd8j4vj+6D
tk4v7CO9ub2v3esToOTA3DGGSVjQQwDBnMudToA5tYjxdsLOeLA2aqzOngkeapoHxLFJxKZJcKgO
fp7WPXpKjTagJadwbW3gUg6M7xg+iHtoNRqM3CJV445d3vVia6jvu4HcWZ3IyQN6uMumuKxELgHt
CQFseSE5A3MmJ42f9pnblDrh6fu6ikg+OJ0e1uuu9sGCRUmLRs1mYzlmb3HyWQoaDA3ON4Ufw5S9
MM1r4C0X0KuEVwNL52JNgZXddPb+SOvRyxKtxd5wl1NzEXAT+FSDaQfQxjWQMwQUDSbl+N6bPT7Z
bjvQm3PAD6zFpZg2YezGozQd1bA8K+PtLildo72mvBaYX5th3js6zCc8xZ01EAQqWx9Ie6s6QGP1
TgP1BFXLnwEHaeBE7OJ+mDOkMLnAKNoHNKbzqziWBkbs/+s15E1rFPcf6XahuMatJLAIVFB0iR3k
+t9i3MCpEmpxeehx9BzI5x063olUtTcITwhYfi3vVZHd7k0fek8TRldXedrGG4nXY6/arDg+ngoQ
ZXy+lwfUOII7vSCziUTG2uEfpxsQ7OI0UKlD73TMXDSCTaQtnHpPEaVVejEvX7AGc5CKg3u3GP49
mX5buxokPMMYp5k8jE85kyqRjcPDb0Pj3Z494EXkBhQ9OGnL+Mai5G3oj40JpZ5aeXpdWehFIMUD
CiyCEAhpAy9wSUGqokaP4H2IGFxO46By8rJiMPtu1BlNew5Tl0l7/V62zAohvyskUAZQjVueBeKu
3UuNYFdrGaQfPXXW4k0om/04QMLOAYQq7br12CGU83DGR1TRTsmV9GdqjZTn86GT0PLJJsim7W3c
5GHg5nTcdKVDEJgqK46HZguvkuu08XqA5OwFWGb1m7nBElYhZg0NJQBWLf3lED21DgVwCc8Rb5Q6
38zVSYDJ4GXq1L8CV84diNXAIdLw1c6/ot/E1R6vhDFlRNKS6IX2mA6rgx4kjRQJNfcHMeKABCgd
lNjir1oUWrvg/33Lg/MwdvImvqr2syu4NW9WQKIW5yvyi6haVMi7qpvtceAVG/kAWqTg5KgMMw4y
AInkjc6047jScpsQ3rZ2dn82tNoTNZGktrPqK3277o6YwhT3R9d0lWYN6mbc/fGSBiHl+uq+BaA2
dGkY3ex2woPh/mWYOw4h2EUegrDfb/ZyMH1/OzGIjInzvul3QsP5KbsdiLc4bdpGigkSKOwLe6gF
sqw/ERT1NiKg1NxAvnJ+Rwkcb3c2QpPUoJkTRtIGXt9zkPBR6ELErjE7HTcN4O/W4JGAyG5ICSM9
eYrKQfcjtIuPoINgE0rCx6tIqVnVvkFK5xEvwrrot/WgtwCJJpdn9zHTrhYqnHpGeW1+FxbBSkgq
R6IggFAPQ1oGb5dnVag5NDY8lcDRBkkcKoGd644EcrIRMxubM5O4rdwnKCGVafKJHrh/TaX1rM3K
jE6TNi6mW4M7Jz31vJrdlCDawP9LS1YNNnRIiEIhK6iu6vvpvekGGLbCHojxEHZwO2Oq6XSAl0FM
SPcUxWqrPdUcsc8MRtbFBd7Z8npvxdgquR8GCre79mrRiqIQGk2EUzRCmKJ2EWQWonvIp1o7udB4
49cXr5jvpsBBI9HwEO1GapJqavSXjI1Eu8b/P88+lVlEHqxQ2lW8ggd6fFpl9jFrOP9u8vS8XWv3
OisCej92vNeinUaH2bewXeydGF+dH9ihfEeSHaA7m8bIwU+kncKEWURoMV7QTXVEpnlYZf/CGhqf
h1+DDrL3lzrLOKrOjYXbL6nXnkqM+JA+tjy935qIpVqOuochFs1tWmtUBLneXTFdPV5LdLmNUKGd
am8DXqC7XIkHN93vMwm8OcARo7Zkrq1FpLx/+peygXMvv8kuvy1Mzqhx6kNNoQgOk4dR0kO2J5+f
fWc8u5YZUQeLVOgxBwh5zKHI1PG5E7GEJ8Pq8Bhkbj6G5JWMDhVhBOKTK4PrT0KINHs/+C20MWMA
abPEUlPMfOjFBKyP51MTFTde+UoPwsKxVD7Lv7/4Mxgh7iDQjbAP+oyHxqkkKEpXf7AgpxSAh71o
ZAABnIs6gJSbxiGARPYdi5a19LW+M+Vu5+J9SG0XyjMqhOKRJYs5gf1NyDd91CytSoo/iJHApbrQ
raEK/qgv/EgRry7b9CiQK1ZxFEhzD5XitVNjwLSGBmNtPCntOivfTgCgVTIJBx74kcmZrp2UZRc2
6dhNnlPeUJZD0IAbmm51Cf9Sam+1wjdWj6CEZPi0Ot43ZxmM5fqYGFxTIIrPPbg+6Wx6PGz4x9Br
pcEl+eIdH+pRmxl89TDZv6HR/8MjAz5677JA1r6JtfoGj7ONThprxCj0b5xR/eLG0Ukm2zCi8+rA
XAoPQ2F3ip8Pmhvtjgd+aEiie4A1ixNaGZZg/UOFW8JxlknNxk9YuyB1Y/p7baDpN4a8SUZ89d61
p/E1jSmV4M3StO3u7S0Ue6QfoedptzLmkh4b3HPNUvxewge20Wdq12Vq0BSlehxoMYYdksP2Xdms
rqSTYldZg5awW85tkY6Bx84Eyhz7RZfaAOZbwum+3JcpRwkvUueTWhg8uz8R9lw7qtIQGjoYK6mT
EO5kHA0G2NzZKewxim4/03REt3yx8zOSG9gjpyzb8pXhvA4Z37EyE4vQpO45cvHQKWkD8B1PJNuH
lKU4AVS0/EOSKUoffRQGXo+w77ooRC42O+oPhpWr+IXmIqgzOQY8VeLccUljnM/XWQb6HLGlcZcL
CFjdxJWNU/UduMdbfeptWvba2lfbIdHXbXXJ1vuLY/S8OdZ1AxGKONPG8cF2jXu0Db+0TLZ+IK1H
W+zaquOlMCALDbI3kN6lyufjs0NEbTjGO67EDYEm9v2lYP1xJRuMl3NV+YPmpQeimOdVhWT8reNC
/V6890kVnsokoESXwqOvHRSCR4Hev/R+xGe0kMMcTNA5le24pKSmOn07BXlCzJhIEBHTl/Z1FDkm
NM//aLdsVbKSwJ6WOAnyEDyXC8evmtm2lJM8XwyBJsNmXRZwuRm27stTJatieYUena5d/nZi9r+/
E6CFsgtUcJ/EshD5YY8VOWpziVXPr9QYwyvSSDSUPpu/y9fwzpSMbymTFA+H10smlD48hkgABbv9
1wrHVSZNrk65nZ7Xhqd7lrOHvpm5b1RvJ5s/8lHdJNzJheKxbwIDe7nhq6OVe/e71B97eEFZLV+z
Vm7SHT21l8wNZpt6QkGVI3Na8DPbdsgIwY1HD/Rqg/90dQmoDCF0ks5fn4l8Vx9f8NeXXU1I8R4q
u4WX1LfenYFq7PnwIV8WISCYyTny94+PfDlwgg38rAjdDvs+nlbzEevv94mYr+4UQy6+iMl6D+E3
ruIBbrQcPHFcL+p4xd49c+TVf297vMcBvpPr0Qhg8psWbh1C9DSQ6JeIO4yeljErp+cjTYM5r75X
RShVxtEREk/2IaipzRY9e2QOYtHwpwYpQnbRFbZCMKc2cTJuoUFqFW/NSVEEcJDhBecntu/sMkXG
CR3RgHVnGey26U0q1ncgoQ21hxS9sD4/BM7kp9EaWcjlbZ+8/B2HTlbsJ2hfrVQfIsXKC+f2EHuP
WQnn9p44dH20ypPac9jqJbgwUajU5OZgCCVxvBp9ghI4Lvqvzw6UPeMVFacNnAvpOJ7vsXm/s0wj
WRdPU6NgpEzHv/dfwcuA9cIfyv1HEnBHPaTb+3AtbbhSJ/rXiNfXl91bGvzk+6rCZ66U01ZoEGiw
hZ/azhOW7OpdWeKxejKOp/KcOh/q4A/lI/pmYB7l5xEOW2QZ9L7F8fyeJcz4ccstCD6zl5aT97It
3+u7I8S8Am1u/KwmrzMVDdES/kBsjw8fjia0pnqp+4CK6yMHD3p2b8Jzwqsx1UayQ24JkdJdIKSr
dIcWWoRj6HCfNsaR7/1IiYsZ2YbW8Q+kZpXDDZSyRfnfH5wXswXap0qR1ccU3M6yV6i8TGvhKQ5p
6LmdzN8rRhgj3pWCKVTSIHc72Je2NH7XMPOjvGg7IoPu/YOkjSTlCByR+mlfIe+wBdnNnPQJiziX
HeryCfi3/YnBP+qbkt2SuLZuP9nJ2DGPqHx/KYPS/Onl+joJIJazd+Y6FlPOuI2XQ3znwvK8PffP
heLMHiJ+AjGFLtpQbgPnTmZiSefqA9zMOJzHf2wPD9y4IjmuGxOdJacOgpPcNzIlmMlFuoBR4doe
Di3pljqfBMTfp5Ie++chndCzylGNou4CorMenvqQQVTp6571gRvGgy1kTu8twOgRaudgdYdmHiYL
WcD+T3RjPv/cri6c+XJ3nE3JmBWnwaHYSMWNNx5A7Gli6MwEBly21JHeqMcoGSetWw7Qx65RajZJ
UPXaG7xgl0gJnlG/6BPWDMpM6pojxySLMVLpzChV7G9TFRs5/Zzd59LXe3Zk/AhcLv6gCf5xnNn2
/CMFWNBskMUzNR9AtL6BZ5R03G0BFD41SXEJL9FEYnaGOUKohIX8KmigVThUnKkU6J3ui+bEiRGo
ZfykdvTNqaA+azomNBf8mF1Y6sN5mk/jWcKPI/ZS2j97ynf2OclcZ+w/pH4CqOTdNBdeKOej3UPT
xQn3kL2txtBRDWUULcDtZnPi7b6Jmg3+WU7PayKoj/ztT27VUmDSQp7O2Ra85FQm0eMMgli4Ffea
/mJpRvQVbCTny2F7OjsaqEoFlDL7Y/Q8IaOY7QP2E4At2m41+oPZG7LkR3Cy61X7tMoEhi/Qt867
kPfduc/nvVyA6UY2S8qwx/FqSuYW9qFyV2wbikmkz/QKS/UqvxknbXG9OUH8wylRKBXxU91Cka99
eeeVKfTqxNWB+H2ze0yH3JTAJEqzc1RD+pKP/h+iAleglQZUlHX1bvYAZc2xBMjr5VFpkQf1RxbR
o96j+Zvjvw702Qq3UQMmJfMvrPQxWJWY6O5FpLe1b27eSDdF0z0aUY2QR3iFPR4X5ka/LJRBQHb2
PcSyTMLsR1q6dBqzCqW/SegAvNJ/g+grUMkNH/qAXQKxi9vDSRgj9c9gkYG8lQI9a6mWHcDd4FTQ
AKH4sMAnb7JSKRwZf0PiLHmOGWwruAXC7bX6cMAm1sKL2QaSSVRBIxbEATfDBEPXcwKKuEswdQCl
+pgj13Lolsh1M96+RhJOmx7FwXOyJDdKduJ1uZ8lVYd/74w3YJu+Ade/AGr2nOD7WBx1VfzZsS2m
2g1n+Ws9fmWvWRTXnEZvfjmAyOVohrmG6CRinYrJvN5AzMvjigSmLcUZ26MoLredoqgPqEROL17v
Obm/UeT66ajf1RQtw9L9GsWMZtIzsTiPx0GBNfVBc/wta22kMndGwXAKVJD9q12YwO442u3knLb1
entVZbYmfKKLCGXzaIAC5I1t5g6bYDfeLMK5weU2n723kkj/pblz5n7DWpX06tRkkLMYnZf2it4J
QFieHEE6DimrMkvEz7ijs2RxmevzsWeIoKUuNYN5lVWQaxs1RwZqtTdAIZ5Uf/vaVA+gM6hwudfE
u1zjWkeWebg2STd6jqt7CmLJ9vN2nxfK35989lv3QCdltGtK8IcwGs5gxbIvzqXdgvDnU8snFpm0
nNJ6elNJtrGpxmEEEfHOxpa1Vvir/o24bYsnyaaz8+xdBjFamSuOab53273oRRdaYaSlEDknULO+
zbQlajFyonSliPRKv4jDCtuWGoYa7uAfMBM8NxuwGZ5i1BCsUWG3R9sklXqzKbHGPMn+rAxhwu1b
vv4GzoFUmApHzCJG2ueXmJXh4sXBs7la/5Olo75HsZp7L62peibuxAZ7colkHOFBPCaKG6Tc2e7Y
G1Pd8FtRWfuoM3vyJtae0ubpF0uUVJiQnQoBqtQ5IX5c8TBKp9Rnvi15Iape/+FST2jcrQ0yPsyp
u6BN/oeIM7ymQzU4AO9QnlsAVUhX9DZx5Q/jkY7IOR3Gmb+85atrjkih3O1JddjzXRR04UNPQkqo
wH3Z2NiMctsJ9qKDk7A/ifv96tUkYzQDvii5o4cHUxu6Gi7891ZQLe04APaMUC/UlkGmrZlFj67u
HsVFXMlzlkknJ7brzTNTfv9MWdc5REtgPUeFLYdtj1RfotGV+Sq+TyLJyuq9xFPiJV8LMMPgTQPz
W+N2XD+tDAO/5X3LllEqaGZITBFQlVZ8+Qza6oTbb/GsVFAmZ/SbLgpbjHw+mhInOgMpwblQGwKQ
Dw69l3ow3Q8HfgJyoA0FHewFvSIla8zxXHRpW94UTzt34kYBM0jemOAbjVZSy+K/ll8t0fzOXUtE
uCkOR+9ePpxF80Js49L5EVnpHmRNt3iNkgKZ/e0SHqQaBHAaB6FXZdLVNwgPfPBXCm0ln/uAoXw+
2KMC7Fyv3nZMQyU31ADptdGD3V6d/Hkv3hSzkNrAm658i+smQqtTW9sZ1x8Ol5LPPnI74Oke2tIJ
0KHVJ38hQNueGf1YPDtsmdfGjryGAgg8i9ouiKxPAoBboDnugbAsze+PnKvtc3TXMeJiPbAmQez2
78K+RMwFsXCc9Huq0B7phtgn99i8oXHC5gZctv/RdvpaOpeQZ0ZsMxObDIvSySVOFPoMcyfOQ87D
TcIx1yVnHivT5hb6iaw1yx081IbjF8B8G+XfOpjR3NaLxgGnm9jNz6EGsTAxHBqk9Ej2fyoRKoI2
P8lGNYvfIPkR38BbDku+m5bXsWrrU8D8f5bKegaVX1HPRmM60s21dewD/zCBJsgR7eOqg/Er7eZa
uym9ZvIdEq950xW5MNg9iszNiJgqWlKDYZtjX2oRakPR+6Y0nWk29v0cG1LrctknCPn81W46UJwN
Irm4BBMZvosk7OUeRkvcEiGvNfQePaXkPWB3Cx+IBWp32zWkdLVM2LvlAb0Te4B6QlM6r2Ygv8M1
Q1N2/QL37HcGf/dG986TaCqb/PNsh40Vh3pqi9lNOdotslly1QjomBtU9S1SGJzFToj/hHmH/p1m
mQzFbbUcgTaiKMS2KaYGz+E7qu4B/n41GlZkqmD5YVBFe9EdqliWYFqrfhNZUYlHNc8naFvfvgPI
tAhmDOeMp0bVXuiNYpnGnlXcYPfLjb5udvLFSgDseLxaTnfHBdUqsmyzPRzVtywDVRso32a7lM5F
ceUBGjsO1dwI89lU7tTgygrwJh4+PjLYSOc3Z7AGFc3v6DXOXnv/pKGYq6U4VWN2EZPzEqrpDZCh
dvKvJ7xiL/QtGOAvmZI71wfZsGVt/fmV/JixkNhoK6PU/AubbouXsyN1rizfnXeIXG1ByyfIUi9P
vQZ9d0mHuFBSYOWfN2T84QkzJfRO+TmKkTxu7EHvt5dRpMaf+Fmrgs4TnEe4TlnRZ2sYUSpBni/E
hU8KoPQOrCbC3J056ID4mjcfxuU//lp0rxGNpNTGMuMEqythSDQ5cdi+BOgWNkFco9jHZyK2GDte
/edbWz+wXYi7K3EL70LquMCa7e9vFpbJmIBbgA3L+I7QzXcbLXlO8yI8UP+QjO+bVd3vk1CCFsP6
Y19TGzlAMpPOgC/iXHuwaGMbJNiud5M0Gaiwf2af0C8+Kc8O3kC2Y6EbC47GHcxWfvDYOWJbrwiH
prJ13xFi2ANRM5nnHEOxuQquwcjdxz6qwhOam2R1szEiJtbCNG6kWUki96wJLUe225u4RuhTgpTV
U0vXqPhJ1MkJN0iOq67G0AsFdU2YDPbHycuXUcy+UV0jn884CAeZEU8GFy6u+kDhrBsh7QpQ0e23
QaAmJH24amfAXNUwy1sGIuV+Eg6H75dtaFl2HbRdk8DauFWlSlT+B3QSxcwp4asoWr3VkZD7JcUV
mwhF8aARFTJrg6YNezZf71j0vbPNynNqpbK0r5vEHgByXTUghy7Fv4bPnSCyWYTxWn/tKVQ/I8FT
i0feyzq+XhqzrInXqcIvF54kTLWf++5iogdzdxNmIxL347qC8JtRFXUIyS/PfOARrh8estgGwMyS
Jp76GkwDUBgc5y96p+Snb7VC87bsLnNazxleDvIciIPrFZyxRtq+hQHwJ1Wom+MtuyhNRvaNEtKG
f1rPtYuvvlwjYRx1B7oeHDSJWgqqRK9ZwuigIjJrqnlk6c3RTPX5Z1FwEjRtAro4WMGcsMzwWp8f
B9cYvuz7hxi2kyv3y9S84zpyfPEi1etLyomOBuP5LFdf3RmtShWB3YyqwFWKHB7774U+1M4Z795Z
T9BjsZHWqO0Tm3HvfnzDaNOeIYbi3Vi8SDVZdy51acI7j9L2qozzwQevU5h8/9w24EPlIS2j6PUG
4vDJTTp/v/M06zmtzAu+ISmZNHbExZWwm85pY11H2z6B5uxRUOp4xH+sMSEcwlmT54hKdYrU9MxO
kMLrxFLy4HLyLj2X5at/7RHlCzdYqyuy48yJEQMX57fBEQLQP91E1sutytiBOGyumw0rfGLk1SBF
ZOZnvLAQ//HIBQS5EZyOQFSC+yYuteppVeByN6R9LjsV606CqWeovWOEUYsaMK0EKRD7OcihFfbS
pH0sq9ywiC/exC74IU/RrfPQaUkIBAsKKlFX82QXm6cTEMXZJwEmbHAw7J9jtKQnyhEV4/tt+lsH
me8nuQgYjNOFMMtmSJPCgc8ZIHy8INiAqRVXunYmgg41ZZimCXqFZI21tdOFznVY4TQTf6F5myN8
jiKHSzFKd3PtSAYZDEpjA/GL3IjIKC8hY68gBhQcf72hgZtPrkyHwlPRxdWrtgYK1w6vgpieDD6g
LmHd8AecOieh3al/cGhAEBfwcF3V0P+kcEjwEkb2w/Re0Zf50oMsgkn6xqQCOTuaKOE528Jl+zav
GTuckM+vLystbyLX9EBZHJhZOAqjXfmA7dNCJWw0QOmyQIIu5xc5CNS5NBHB6mu3hSc87WAS+UE2
S9xgYN1oFFpmSvygl92QF22jnRL78j0c8gBLt5sUkQYVoVwYB17JlKCotE0GahtKQuAdIUoEU7SI
ktUWtex1qXMJChUrXYctXBvh1A8WlNRvWtmhrS7cPXa6UKSTAcbvPIOwLLdrwPxyJPvbake5eeXR
ZyTLn9doToQL3a1ORZZNrEpa7oC+yr2G7CXefUCVQjneon+P7SzCKsGtN/ijS5FC4mxfnN4cOvJl
CzR0QoF6a90jt/PvnK5f6/gShuyqXmagf4zyKF4g/8phHsP6AQYahB7eX1MeaMvW3xQQ145+2knb
vqXiCwX2O1DOU5YeBQBTEy5XP6xdr4PJ7j0gmmOPFnPNf/iWMiGlpvdaSPdC0GA/gdXA4UrBmizR
kfaaSBPBHnJcceu/nQU+EO0XAZ2cDGOF8h01R4ArZW5DVFOg02zTNfjFkZOgtAz48nK+FXIJsG0S
K51QsfdkUfD99lpIWVWs61j2KVcNrtcxH9roFOCnAK8B5HId0PdtTkLBv/RChJUx+4D/tTjF3r/m
dV3DzCxb0UHAFD+viOOevWs9nSmJLPZLxi9J7JR8llBPkiLi4sbOWTrRR+F/wdNPLLUKQJkW/nB2
6AvNGq2P4ZLPXOScD8u6Gg96xFkx3jTP+i76aakgfbNn3uWCtVQ6Bj46KJTbl7Yw6AlnMsS3g8AP
QVo7GQmBN/T68Kj27H4WOn0ybc4TOYiuwlRMaJHm2D0uhIDNc5cUfWLncLxw5bDgyQh3nQoCMaVV
fgWKtOw0CTKU0UJYMF2K7r4YhuDnDEtmW5kqzngd4zyF1GOzelTizWYhaSgFYyw0VL/SLs34plCf
GvYqOigCVhLQb0jqhb7avJITi//q7zTL5cKty51GdSRAe2lq2XC4D+zGY1oapn4cxosHyX4R9/SJ
uUulz5LtM1duZBcc4P/FoPUUkJVb4gWemMTBhS6oDSb4RNbK9BM32NO/Uq+uDXfIaq9CFWbD1l1p
WQK6E0SZZDkNT39V1NIb43y70oxSYJtPP9Y3asczsCq8y2sNIND+MX+hhz4EO+Jz+oZZFeyb4Eyo
mfsYhuU9zF9Sit8PSi10/bTkhXoOkzu+dJjaW7+T1BT+porS2JzFRxG42NZdtSFk5O2053WD0uaL
JtGdHHooIizh8CtNHtc3GFlnwt4I7WW6vo3kziJUXRyQVn7d4ud5P40lrj2Mc5owTRVv8lBi5dbw
Qv0ahhvCCZ8UmPoS2p6jYByndiN/h+dtlCvLHR1Aj4JrosX10Xxc7A6UdDhvpfddkT4//mYVOuom
/Wp/tBlLXqYPaiKKme4Yd+teTsQ3la0LoL8zdffy75TKiEmv0eBoFXpFQYCnf0fKujSJ+bhVw/kJ
nBThDj6PdJ3ocWR7gJz2qEsGMWBF4ZSVMMiRt6jTS32j6fauTlEAp0CfUAc/L9U1Jp7CijVJJSiQ
V+Ad6eNvMSFIqFEDCMEbC69EIui+8b7jcY3xv7/0HQv7v+eczcaUP0hmsr/35HyiT3/S+CAluerc
TXtNZzGk70oaWHX5pgOvDqwRy1UV4+5vqnXtJo3+j2yjcCbx/2XLMMFvadQOfJ7mbWsklMVpmK6N
ne0QBq/Hl5zhiNan3tec+wZ93nMEy/W+Lz4/aeXtWQMUIhylMde8dF/pkMr5OgT0qbVr7igqKH0J
w4RA/jp60VoavskFO8FdTJYtVQB2+fjHeoBKpaiAR49NEMjJCtQM3TIU4AdCOWeC1k7lr3gmkbMi
tf8UfLt6W8qR1WCpQLpTZXD0ltgTTkbLhigMLFEQRBqWAtDmCts9qLADKPClUgNCkWkv1k3JKdJ4
+olrP3rV4d32icpAmlZk7xCe+cManx5VkU7DfCtUIE2QpvbBKMl80qHz4OOgwf/u56Xi+sePE40p
HDQMeQmGRCbUGQEeOMr5ny4UcGSdjokbElbSsEAjInaKXyWLTbE/AKqfcy6mv/snmBPDK/JDVzHn
6rdaZHWZiP9FrQxmVYXYDdpXG4cnV4TjpDsjKRs5RdwzuOrCZY8aDbYGL3eA6PejkQw/Hp0J7laC
rl2o34MtcNiZ4ToD33joPGWH+HTv3JF7geOSJTGWa+bI3Si5YBDo4692W3w80ZsaONqpM2rrY/lh
PCxvw/3Ms/Kf+QZSP0anI+Wnpig3u15+iBmMnn41RQ4nFj+N6/HXcHgfN97IkxxnXz6y/gWDvDSW
57LOw18DZlQ+IgYDGs5h9QdEaFKJ4BhLR9sq0s0eWpOkvxgyAjqwOwyFUn5fxwx/Qlr6cZEun//c
kz7f8Nig4tRpXUoAkceXUeP7+hS99Y+yBFuGwBAVPEw4P3BG7JPjw7fnu5BYTV4rC1U/f7a6Rki9
+Lmo7iolOTQF3tWLyKfUBJATk80UA1ctUfVLdvy/ZSnxZuurU+xMo7A88kVeYt1TzVzm/rMXe1NA
TsdCU3OBTTHMRAehtSfE8VGpkQTFogtgvhH42kLffBjdNAexVfnUSDtU4g1n0qWnxAa11lKPImfg
xno06GO0OPbrIZq8LdOGf8ZRB1XP5VfGbo0Jz/iyFc+r7WqnjKRySFITP51FjXFEp6VPDiD7k6R2
LyyWOSwSBklTVeOsKZ8tTIpLo5tR/9s27xTisiLIWOSYnzD57OkDhaFiDJbzG6Zp9Ff5j6EP5f3c
YTq3tgsycnm2GczmqlNuvJmn2pfcEe9f2lvGI5zc74ItDHGwDnzzPBQQuX8djyCaobMv1kYxL1Gr
Dr2oXC/tfhfLRlPgd2jIOJ3IuGUMhtCsmhOBGAPCohD0Enz6Zv9HF8ilHmHfsEaEqZiXS10qyqeB
CwydTLcnXPQHZR+iLtEjEccSyk22XaDwZWPfB9/52LZyeU+NCG73plxVHhnw6rQvxFGIN72YBvHo
1jlpPM3lCgme57E5yWjEwlDJU5ZZVRCI7/iLyXyrqJGSZ21I0+1U3/uPLi6LR3j5mWpSwtELA18u
yHD2i5LgYzyXUrTluUaVQ8g6ySVwv9umGwkNHIdErDLLFmVzNvT6miR9UTblRxrb8kmaqdPVfRhY
kKXGUG8iejs6SDsR65vMNOo5UnrgfYMz1DaifT6itPh68mCXSR/qws7v14O2bSWdMlHDuh3b4jNN
ScCh35JaEb0WWg8ntO51i3naFeqCPJ0yu2XTCnfgsRfTjDAHyCUxUSR+ZxVc5C6j6yBjjkGbfBxE
GNhCK5O14xl62qQINA4f3cnZy+W+OS+9AgFsnsdRT9xhpnwuMpM+LPh1RPyBtmG1pLLofAPvJsDV
bxItuuvylZrVrPoYYefFi1KvVI2lvbI4dtxW5oZAc35hmawE81hq+pzl3DhPsws19FL0sPTGD9jc
O5dlumHrT0Y6Zt5fdMcsmko8Xyy/X6/esB8p9jMvqJh3gKDFYt9xUiCLx9uPdm2XA7XBKCU6h1Yd
VhJ62oas03xWIxwOSmsf4cIxG/FbkcsBkLLejA/dFirTU1ZIUGOiAo23c2m2gbQk8ipnqI2aspkD
VK4/L0m1awUQqlka5/8BbGVF1InieuaH/SEKlnOgHyHKczz5hgXzOQIhdiT9UExnBdnIupLqCR4U
jZYDot2H9zMuU5BP314HvkPJX0+7yz+vbWHSL6U8SGll/0IoqybJM8pUGo+l/+Pj/quv5qutZgw8
Eta+JlEHLYz20i2oxhM/OS1Cy6hM9itpOBtM22uACY6ZrrmQElTTfRBSGAXqe3pf7o8PUdmeib7q
0Uof1MwGqL399iukCiy9qgbyA4oToSzei7gCsSLafL5imqCHgX+L0XMk5n+zFPDP6dLU66f8vI0K
n/CtHXlav4AJjlZ0GCkNefuy71Gqp2ENRokqUjSPbIc9RURxJrHNq+oejPvdiEchbv/0dWeawOoq
2416e1BNqJ7+dvJQogt8oQZn22BHX3oq5weAucGIb3wS0gukosWIKyQIAtNY/6bPdCxHSzNd1lVI
wPMm2w0pNOKUyOLvszEk5B3ba2y05jFyNkAgseqvTboy9nzFD3dWTTvPVd/iqedS4xESuRghqJhl
AGxvHQsLPw5Dyi5MkCBiSH52uJXcp2BSvnzLU0SF3JwOd+Hv82Gwv3pYPGZwQMc9vD1QfPsyaroX
F/hPxSxcuuCcVqmeL3dOgTZc9C2mfd3JDnSsHaOf2xW/oMjMpLJXHJD0+UJ+DyN+KwSVS8s1Q0xT
dYT8XEypuzE4jDH4lu56C9w2hZc/dmIKSm+rsDKXMAgshx9ZCkAPe/lDOmnpq4FFa0GvrU09Rx0y
sXbh9nEEGHtIVwOUBEKf5K8i/VsyUyqwV1c3Z4I5go4bgivpWgzNKU4kPzWewbClOgCVlM/kB1Wc
19sch0+hp9FOifZD1ZjtiIax0vFZ/lw3gW4eC/ZcvUSJ/PGPMw6VRZ40QM88dtSNxlQxJPb0XNPb
1ckOzjmQ+s2QI5hOK3TSxobwH2m9zyEEVsFb8dZA8LI9NN+bH2o2EG9F7Enljr45ALJ4yqZf33mQ
ViFH0dr4b34F438iiWeHjRcwG8LInPwawZF3cbNkn1ApI/jMQFF/du1mrxWZ4+qaDzBP0zAHnfgc
2AD8XPejM0xHJTta8mw+0EjQHipaO6LivsLz8yJ9ZW4uOw/kFY3dK7XDNFRbW67bk0whqd87KFMs
Lk0F9AcMljYtv5nT+RUb+X/H3Ml3NlF07DFPKeNgfcdoIgb0x1FY3ixgy2l1VbFKViirQwkPFfyi
oo3nBrZng3Va1PQNm8qgn6F3c0JKNlzKRoDXbakwC7z8i/vPTKxO1e+1YR6vnRFFCZ7ENJeRKcyU
UagsNY7ZMolDn5KV60wP8RUyVvbTvYyHVHuevcr5wCB0oYz8RqSybLxiGAgz1VYPCeBnI/DsYUiA
Hfdj1anagRH344ZEB+qOHKmwOkBUbwg1b/nozc9c33VNQaF17JNnI/g6KeoAwiSHQY5hKxu7hjO+
ko3cxFb9DWOzi1CIhaalgk95cpR7KDkpQjC6vpTZpgPxDmMHGdMx3Q18AFk7gNE2pKtq9yUb5p8w
+zwbH0YbzSjd6ny2Vq28T4qm99K8skav31zHtz6F7c34xiDKSxTGK8hypImebPhh0RSBhFe0UDkC
N8P5qoWWM1WCYsboQHYCYlwbm4ZV0YhtNMG8gDXA13+JokvSaH6nz+5QMvzAXpLc/TXxFP6qPvFL
Saw56q10q6TE0cxock5gJRZqjIeqjnm/R3lvJFRxZZEI20O2d0BS3BakOdThOOV+2M2cT1doe7AO
WhGSn57BkSErTB3LQgnBbG5z0bsdgmhsuFj/RAcPiYoB7YBpFTYup68oPzVfhypmm267FLfYP/Uh
DU5WL5rn5R/8dllQ/dI022DO/2Tv6M7FMzyu3/KcFUkChOjhVLC6iEQhohpn1EbXABpmwMR3/AfO
fyokf1MzJfvzD8SJbDUcimpIzzb5dlRxjztb5sJsyAgbDHLm1bEYj/z4eMhQ/8uSxwatTwLUGng7
TeAWMnOrWTQ3NATRWZid0Vw+F9bxBsWXWgvY/YrW1soLIQZ/lMCWDxl0ZY3PAShtJVpPjfL5QBl+
eO9rnrm0IH5Qqzji7RvczFDEJIuQ9Z6w0F93w5oj8miNewamnHBLHKTPvrfbdeRiuQlTJzeIjsCl
a6OvXUcaGXOsT4JOu7bUS3zn+CIQC230dnPqEGew/pawM2NKaglXcqwfltySHdO6R+OdJ3xBXXri
gGOmLmsDRed80hbDm/u1wzPg40p0jgh/GHqgePkesnWihTGmA24y8KoMel5kbZw6LAndOEORdUAI
Bi0Wyu6F2wkP3Oqr7MFmOGQa2TlTOszkwhUptNuBuLR+v+9A6A9PN0Dr102509NN6BNp7EieBVxn
m4HUS2jmuiTKcitD0EE7KoaEghYxAY0Zvifq2sx8Mb5ToBGemfHkRPJxocKiVckRNYvxwhuKO88q
jJrUwTyyiQ0wiviXkm8KPwdTeL9fT9cwHIKs0h8iMqHIZgL3rbAYsAY9KrpmlN8XT4TB5YprTiSb
9dNN2PHDifUIMZFE7WZwOMFLS99aaBL00b8LVHm/M8TrkM2dhnlPJFmxpzX7W9BFYVr8TEqqy+fl
EYl7007+WSYycofOfGdA3u00zu/gUuDq0R8q/wVnFCQXlaoWtDWC5EcF1ltb5UG9or2Ath3bSI8c
1owlO1ESA+vwur2FxiTsn7ND3wUD9GvJFK5ktEM42olf9kAdogQTMxHqbBIRckAdyo08csqS3igU
s/6w7igAa0iF+FVhS2MwM8KMo5OEQOXjtb08dCbj6wsLznSCgBDYNt0PJKveVugrsmryCkBRWWqL
FjDZgyeNlTOgInXnU+CUY+xHBlERBlrqPdH51siWpDj3SnCRr4NWee6plzBNVI8YycYIut/2+Xkf
Hp6gCPWUAvtNzJNn+FrfyrBn9iORukwByIPltWA9ifqZnj9IlzWESPrbuRqJYV/d1jaPwCTOmvO0
blUzcIwwaVTCCTwGJP9g4S6V0ZUIQm2Tsuhirr+KTzej96jYv5QJ1RvRAAesRGv93F5KAUMosufy
1AZU7EfzhhdTPpuOLs9ofbMH6G5EESORHR6BcTSmpEBDl+oGJEkND3UvfBhPo+YO73EqOcJh0S6i
Xq1I5InGV2vYvgFtSDGJAZZQALJ/0LChxehlERrcTFfLG6egImfCCBSQ1PIaE3DgTlkjX5wrpEb+
G6nhr/HkBhCGaNmbkq1FgfzccC3PX5gJUuGd8EBCzg0gxa48wf09Or537FOMPm2za9XPqzwbdF3u
AoCbZLz1VuCDe1QdMNcLtZ7kfPpWefY/DUQ/AwXjJNKDMQzCgiMsttqwQujdCd8Al/Qw2WXJKqVg
HPUqfFGC0xojMlPhVR74klZNzLjwIDso2giEhpHwauu1YXeN0I08UPozIMWxPIEqrdaZ7Q8FEh0N
ZJ7rwQISntN7E68i+GPE21tcU0I/Lq5fPJnrIifKJ01ix6UxfVRwB6x0zUKYbROhE01Bq5qPaGB2
ifAItAGqW+U6ep4iV7+qSsPsfFya0Qn93RuC5XZllwrtuMWrlmbHyE6Z/yQkuCHjouoGJ5tAIyr4
JRcB8mQMrpl6gGEB/b3l+DOIEA76FmnmQ1LU5FeVH0Cmozs9lgjQgxWHz8QYXfW6M3/W9YwMewg/
UzRUzsQw42FVK3aV2SyHK7yiru/Z8qoS5s4jsO1Kk6JMz6v8zlTV6EgmPWzZWPl0U7wSniG0H7Jg
lRRIFjFkpjKY6lbe9cDstU+mFqMpIEUQxRqk2qvhwR5+sXQ0PWHrOPNMYIO+T2JTMuFHAozbEdyo
tXV3IFrgPluwRjK6WMQrUeTsryF4fYqQ+QoU2vUYwWTeXozrvmGOnhNGi9qdJbUemmxmDMkhyFT+
w8hCyZgPEqzoOlF4YtGpnhEV7dOcpKV3LfwILlA0YPp2quzDM0C9W5/41LLGe4T6v6sXhRsNr6rn
VZzUlq42xYnfeDH8K7g9MqDlICsnou2SamFWjO8tZOL/L1i/yf/i9BMblF6KaND5CBHjhloduGqu
g67l6qAR6TZTU7NEDqtg1vlsRrWBa4DqtzS52P2paIg5DnFbpqSKCuNaNU2BTAU8hOYTf9PQfMVr
gB0LAvL+K2f6X5YP34NjkFUSGdztIYUWkWqP1PztCWriGa+ApantMIKmWEnLjMMIhciauoIrMO/D
3MG6ZyKTODXjX5+rUcykCrEsDOyekc+xTfl63K/5YcH2ChzMaX5NFTiB+Ru4xvn1EPCwxMNFS72s
EkUvBO0Dn4whKHRs+4i9wnXSBUugoNeYj5AQj4huRdLYw4JoZLZVx8jac4VH+m0GEEQw87sy2sz5
PECQzDsa88UnU7zPgZ9B9FNJM7lgQ69/R2UV0XP5ip2QJMxlB56ViwkExV0WdQFE6AiEf0Qy16v3
dLvKoKGPTi4heLhnUiuBTyBK4fmayR5DwZlXHUB7k8thvR8eEjtlNxtTb5mgPwBHXIcmt2bm7/lk
3zwViSI23oPq//W3TBuuYbDrFWlV2dVIGTdYVPN4rP2OTa6vHwyp3GwfM8JDFXabLdcvTkVxpsLi
Ht1FNajuQ+K/IzdSBVzmLbPNsdnWPdluNDrMpSa9EXfc1bcSa+YN8F5/5G4KR22ddq8nUVm6uosL
fmK21nky43o5huGEQsWTbDOd9vnWJn3TIYVZUtXU8xL2CUykiuPqugg8fF7Yx7Gq1esTAX/IPajX
d3HjW9AxCEsg2GBnzcn5wrI98AxSne9Wy1HWDYF9uH09FGtrNvJrhR4gZq46uQkIZb/rqNKCKX1F
iFS1+9o3wm1KNmIvbm2k1hfTGe7DPCiktuiiqvingD3EycRS4J8VkVh9qsGI7DiURcT5sxwddiM6
C5xP5ks4ISNZrgGrSPTDA4Ii9cIjMSpy2iyPnD1xH1aJz4rfCGZ1RO+K9G10lnB3x7MGvhgFMkT1
ISl92PzsK5aoBV2NSCX4XOESIKepJsHq52qvOp9RskjzuFhGCLQsJ1QM5dzdIefAakQzMzfRcJ58
XtrcVoHaECAvh8nQXtNWCGJgNaszTI7aLNnWc1CyshzCRDYgvSByUSU7kqqMTNAueuC+/IFvNPK8
oI/H+Asx/sQ4WqGexwiQs7SQFxTsie9xrxRxyDZefI9OTtC6FOqWGbVSKO+XiI9nIXhUAKj1OjZo
lMXSXDTW2pa9DWJxLEq8TAwy4XPzXiKN0Rv4jmFu/Xm9YyNF2ybE0cchakP2d2P9ox1h7TwQXPxz
ShCGFS7mXKmp/N3epr6l0FWfq6EuMeqxoYP7tnkhNz1ITRhxRPz84w3hpp+vTAd46uGATozuIkDa
u2wVuSvFkFTTVKWhsumcvVQoIU/Kdz45PWdDtfJTZoZkqb/oTz4p3ugcQCKaPhQpefr9/vzQScKx
0NdbucYR3px2c1+gTFwYbgZJa7cH0ZwmWZ2PaHINHtv+9i8JnrNg/0qQHd77AZtpG69M1W6kqui/
uLDVhHu0s//6+okIkY10xUHIoLxBW3SraakwkMv/ucheJfm2bqII6URBXyRAlMJ8L7K+791482or
vr+/4UlCBr4slEwhOCXUfD6+Xb7bgynxMNsjU6+/W0yFoS4AOirX0a+MFs/ySRRZHFJfdmR3o6gk
vMFGC2Ug84AulQR4tzdXUsU6zpBUyaXyhW4zgWnVBcXTw9IBEgptFbUEXxyS54lJB+vsmf0wmUa6
3YXHtBGs+R/MzLngWyK9cf58KtyEVdkfT7Stm67fk8cW2QE7RCdO+Yc0WdFOMbiAEdnu9Mr6w0Ag
QqPCNiRz7ougVUhOZkNRYjXFASWBcJRC+opFK61CzAtfnFdx4+Gy592zZEhByirGdklOs3ug5gMw
oaig+hlcI4Gf6A4dfyofhDCjmrKjHvopDkrbTufmYzdDDr4Q/3IRLb7NOrkbwcgCW+SzOx/aItPO
YTPxZtG2GE4/lbqlG98K3WWfqGm4IiWQLwvoQ+lhqGrDQVat4Y+KrOnUDZBGPkbmmhDGovsFZb3x
bANMQso5yygw8yKo/IV9nWX8tFKLRs78/5nzdEAxfZIrNjksqnQ1xbEs9ZBKYo0KsHs2MG+b72fs
gNr+lylnlYwtGZeuacFZ2J+E86T63gaxeaK+/so9eXBeBqV42PJTYKDL0rCAcMfWezJ1qbK4z0zA
dTqD61aeDkaqv0Ye4tjwK2jCPv6dFq7qZ+TpAYsGkUhEmIfOVjP19ENXKXccYzvTfWD1vtFeHRNI
MLQjvIq0jo91QapGu1akr5dO2vGlefSaQ4FQ5/Hz9rtiak1QbfGI80DbeWF41R2dbnJjG8YVBFFT
bAaNRky4fzBl4MQn3bStcxPlitekgIRUykMnBOKvfyHxnwX4z3Q79zdI6tqEzVDdOYFQGwHce9Lc
mVHG+JVKh+eC02xFlfLhZLhX6UbvbdLuy+Tke0JOP9q1bF/JXfIH3lXQ2l4WFWOEsTzvOyrs/ucW
BaLUYnJtUO7l7oU0WgrEKzegtVqYem7uDFd1duJunigfCPyMhJ6bNPifK06dhnnOVQlYupnF9jzF
xs2wJReysyneyp0gzC7Vp+uZJknyUUu7CHopVdpoFAjvwBOjh8jZa5U5xCqSkEXf3vEZleMvYZlv
gRS/RNTnx7D2clWKRfhERHQahQUIO00CjTfDC+UctjhaJm9aZrS64oJ8/JQWoMsgp83oHXkfVx9V
x6F7lsEEcoSWb/9g6Fn9waQqpMdbaDL0LPVi2TbUCY4zIXYcQoh32+BhNx+MZR+t2jkcTDa3x64S
SQ70/JVBVFIk6IwPzIoKmt8Svc2KcdLd7ZYgh2rEN1/B76kIiwciRjIsouUf0qSKOAMS058hFdxn
EhR+2rkp4XLuD0UI8c5xXMrZmBaD9gLFk+iKRX9xKPlosUC/6HqkVRi7UN2PXOHaJ2k/B1SVctN2
mn5VSU+hUhAUtBiMXhEkkEYGNY4ZIfsJA+Y919vEAF/3UnezkzO4g4GTzH01J/EsK60rGhKguwbU
R62wFX9EhFAoUHZuF2hHZeLDDr8Uxv3aMuJXMzBvf8MOEPjUrRHKQr9lOU+8Xb2GzkBNOozGk4VZ
dx9aEiOQWELtD7PcV6Hu4GJTGjc6PbsXPM0X/6TPUQiZ/A2+eOlF8J+t8khZZ7a9ZXw84EUEZKhI
s1SdYLaGJRPcDIvx3bc/3fT3SlxG3FVTnJX9FK7ZayOSwOpdlPH+pecRLNp2R+SjctVjHZBOGwp+
nAp+v6VFIPP3eRFEMbrxaHIjKh51Nv9tdb6G/QoSL/aSEnCIjhXoxypidnIhNBZQ82SGFwrP7/nQ
phm61No4tA4URJrCyK+FFC+G4yJUnwT2I/+L3j590EIIsKf1PahZ9SuSj0nRWBPw8wTuMBRotRmO
7dV+pfQOic8T/CfKgzdauwy4iIBgW2FctpQa7TNg659YXtHEu1Eex62iM2o1ftbciBxk4VAwQpFA
NSxZIn6za//Ns4ZAmBG5ZEF2ppe7o9T46Snp2VMIdxA2XZkMMAhNqDXfoiLaQpdHFr6vGZU/ghzq
tVXWV+VTENv/qb889bGBKQ0Dvu3DYY3I9l5QjsGHuFzjRF6YNbtLCAul3YxRJ+nIBYqg47PjuUcD
16+dMjDlqIEqwYSYIVuQQR6uh6hpF55A8dc908I8vdoEWsdN+49UggI2X8ijqAP50xZALMUCZBEb
UL2a4jtcZLrRo6DONJP/QPXXjDU/OSxrliYIuuJ+XxCUyW+9X6ifV8P/WqPFrN5Rfqq2lRHGcvyK
Hx5dgMGYm8PZI9RtEuAPllIKImGsve6yyz5cim9h30ZXsqE+rKIbdSLKeIVO4UaE1RkzQ+VREut4
QY/6aNyR3oS7if8mkd6XsicOkVaJzrJINNBYmw9dy+ipLSqp0Twf1Y+aYxzi+Lg+s72bY7wGp4U/
5ody9hROb3PSyuzH0APfvXFX9+MUb3lGwb+/9fLtOprUmzfAkGjF9yKv71G97FXJaY4TTPz/PJJT
ZfYLT9n07pvIF2QXs1b620R+vxYdvZcf13mzQLaD0c5Ri2/bslhGfdrulsggIZ1rVg7qurpGQglj
1axvOFTzdeFotPI45tIf+zVBs15OKCF4DSUvRGoJwrHs0okxz/gLQJEuL1kxyepsx8W6S4N5VDc+
d3c6Wl97CMl8M6IkOeZ9X+FB5s/uPfvOvoqA5PulgySlSkf25VJPSG9RF2nIdEf5GenZt5Hl8izW
YdAazCmHEE7KIlnt0R3SXTRZTa90H7cRzwj+MajEpfQP1lGstk6w+5tMFcv0mhypzQaNgXQIbJWf
ihvPkrisk2WxUr+ildxf0p1ZYux0ttIKUJUm5vvxmxgRaYcqol2ThmwMpzPhy1+SwjY0LLCI/+QC
xIMRv3TKaovD8NZRgH8pLJ5XK1Ohft4oJjORjjMJ6xIYXeZoFwVszRFILIA9FFmPdxp2Znqu5jat
nQTdMTcHMp9MKMkCOdAR+MMky3Vax1dUyLx2dwfT9bL+mOUeRW928t4VKIz3dxvZHu8ynYLReP4A
kZO0m6efDcNp16NmU03Tm+Nq6Jl5COoWlLbCAMRE2yVI/aJCrCpTCNj60kLK1QwrSVmDU2fO27Dy
b37//5pfHbbGuHXmQkIPzieHV/icKaZ5uHgzSsJXHE4tFT4xDuQhMMhRztaLFftDQDm3gyNQRijJ
uOUwZ/PjoNN7IGknbmXeiVKpk9BGGcHA9JBb4I1cUlC3t18tPQkUs274I4+dJXlOd3YcwYzYlFpU
jQgQgrz63BwkMNoL8UUTxcXa5egIBKJlvDBxpPQT1RfRO8p6QrGo9kBbi7a30doYkPeLwVAItDcE
bydOM8BjP+TywMUmtoMZQkyGyHTkg3u/0axTNLz0uUQL+A8LwhVKe1eUybAgVDPxNm9kLHsWpsKU
pglx/PF+qztBRrDJ5yLJ+8E7yE83vrDBp2WNRdQNJ2pBlIfeqRluGIov5FhLcbzh3H+mHDNCR5eI
LQx39ptw6Kl20SVgIGgpqr6T3sNhYu2JLEbSYbS8K7PKsJe+x1L61aTVmsXYTAkOz8MP941ZpUBn
TiLYHmtLP7NHfZeZtiavG/AdJl8PgQQtnfIu4Y20wDtVAYS8G1QaCUzJk9RvbT6y/p16IM8jU0MC
5ANLaesxHIj2b481FMCQMCkadGS8ITzRJIVPfBwZeehYh0xm60F1545ROMqV6FFjLbon0iVzQ7ug
Y0bLJYLpsC7nRMulebWCNVCFD52Y9DV59to5rhesqW+bHIsSSnsqJEqIW/5lGdELl2lRFB9NTz+r
q0m1ZX5J4Z4RZbNCKr9SwvBllXtmR4xfQS9cP21MrG3rpplvZbr0F6SkrGSQFxdrx683MWk4C20i
k4LktyA0cp3hwhWamq2ntkHUgcm6bX+dLITfIaP6ERIAFTAVgeT0UacZejAXkqxGviCganKhoG2d
Ft0Fk54iH4hoDMF5jKZb1ygo3wpYoXwt+xaZkGpQQCsaXHou6D64FB/UbAaijT1xEo+WgVzXbdcW
tUs9jpIaTaW0JHklX/EYki89jIUd8LRPKmCQDYOe3856AenlRpbxKYgHbMT1PbE8MrKPra7pnopd
EaDtdzBPDBXPtwQNzVy1f2MPLy0lDc2xUhXLCc9O7MD0Q+XNiBogPScRaKcSLWxv74N3xcW5U14c
kHQPYeO0CO7911pWTVmrwQ0q2uAqJv3+93Pictzr5UnwGM5/JMnAf2nGNHqvnmU2JBTDtH0OwOgO
7NKa+hO8V97FszJrMYRliMPAC/jl99/T20NehaZ+tdG9ayLWnuDdp0TkO0qrPfBklZLZTKF/hHRQ
4w07pLJKDIfqE35iB4OBM0ARRpnF6X42ezfs85NEYvCDeOYAdwWOjH8N8zqr5srGy8FQLJyT9yCc
RSRvNH7bAWiJVd5CO4bL9+JeqBiqLSUFzH0ygqXmzLV8h7cZDEixrhixUZ7DmZGy4oRFwzIVGHYb
jYDMFgTyyP9K4CvliYeza8+eI6cm0smPZBLP3NQofj0tONbLjGkfzfntx8YoMWVPyqxuZSf5dqlY
CTZxXM/iwdz/cJu9x7m3/qfXjwzxwiDVdlXAGSesjyifSNpyeXcJ47m9zGPgGzSQDEUg77gTrB8L
2UeCUG/Vp8rxOCayhEYLF7OOEyP0A70Tzj5QQxDFmYxDCscG2evDIPbZ5KNCOeDfl43BHoSnSzKy
zayFS9UtCcgXXAveTStR0ckDzHHNdceFEPhhy8ZvSGbyo1QaFtIOKvHXq/IYFS6vktOvMwV2nQ4f
XZT9JmwXkjLZO5vVg2QgDMF8DAiYawnFT7W7zfx49FkC/CyrvTv5jBg0SfHDbna1324BJ0wkH2+n
GZOerOl7ZdMv8K/4pIlUMfgUCY52xQ/8gOCDlmwC9L5/Rcpqw/TIozjkkpVLpTZAn15xuK3vQGIv
8792hL4CoQQTsuzKIBGQRYycs8+M4nn3mhcGHrVcBcAMMIYdDpwzS8GUlqx3caKcWDDoyJ6FADlF
Il5VUJZ6YgC7wHIxIx9HQX/6G/RIpucqeODucAoXls0/Gm4EMYO0sWz1cl4owk9gQInl1H5f9Ajw
i4WEHdgDJ9RjZfL+i79qJbad3yx5tNcgzMX/T2Kw8WdMRm4U011L8GuxLG4zBTOA0lWCTEnzh/HK
UVDLa4XH5v12l/rx8vEwi3eyM3UsseUam1kqvgU9crTJUz2TJJjgEeui/i/yDQDhSr2aQAQrx0lB
AoZG+iFACRevphmpb84fEdd19P3pCwnCfOvPzKz2tTIH2B6+UsypbTW+YqIBoQTd7V2JLFnaisZV
yfWfseG/IX+A1NKjaL2FU6fvb/VrTRFtC3rRE7pM5MMl6cu1WdE1U5WjQ64rB+06REmQnRu5Dkcr
oQIK2C30YNGBNvIL6kzTu+OvhaV0Kkbcl0PaeTyuWdHqRLxy1aZAbosHAoOfVDjkSYfgZ6lNlBS/
WSQPbAN4eZZMojr/Nc9+zPOhamrI8kkDt0qh5FEW1WneQMcWqu1Ra0rpZ/GBGzVASALCLTNlcQ9p
2AJcwLhTEanQ4K8GTEs4/zNHzm6hrtUKVrAzariHRjJNoEjo0asJMOxVPrcVN6Cv3mPY70vVKxlV
9w/qrO/IIZDWMgrDOSJ+h3K80xPK4a1OfKKicFwx4yic85v2E6HofI86zxeq3BVQ4CXX5OR2cAvW
2K08HJVjyy+8qBPQVhBhhlAO5KSNeoxluOICOlM0ve8cIzCUGm4wURehDlzkFlIWAEUlIVdoxrIU
XKnewXfHUSnJj0eaclRH9DBJs2h8BBAc2czkV3alwVSrcu2q/PJGmtU0Pa5AelD0gyPMbpzoJ/ei
v96px/gOFkaAa7kOgk8/CFcZq+IAjB2+cY5r90q3o4iMoDi2VgiNQjDs8MnUeh+T7O4vi9sk+iO1
9U4SRJrHwmRff5FYy2toqixKL8eo7AOFco5dHCJ0gyNyXrtfeDNloDPyqRVH+t/aAZUZCQGL9ap4
SX9Pakia55UAdX3gdnMJBHcv4mycxa1dKFbvwNlXZKPpD2TxCMk1mrI9jd5oM2EgleAyZxylB+1s
4565hNwPM2HvPGD/UrjBTF6Qxj14tW1jGHFf0gLCaM55Qj1hBLsKwpf61own8roC+4PZfOYa1Hj9
E0V8jW2wPHURvxJr2d3e8wxp34DiC6vWo/WatC4mOog4kg+NC+K5svHXboC20Vhi9OrIBpBvQhZE
MI1z6BPSbKpGUIbzG4CueYLNVhB/Zb+WMKjHyUbeg5lyZnp3XA2JD6RCWrdBrFqCpyMsS7l/w58g
zlsxkLjdfUk+J4I7DcD1jF0RLlSH5VhMiHz1pRIUWJ2vEhqPxYOigl2hvzStlu0HPahIK3A0xhST
u/Lk+0qUN3qKSCv2Ka6FwexBNTaBCDrG7KraEjOjJ4cCsAP2AdHDPsKnw6LiS23rrer4TcmDPE8M
O7yI8ylfkpee/w+jjjdx9Q7uZfbwY54U04W2xwSpAPHVJdxUHQlT42AWrHC/j9vfGwL2nG2bwDvE
gpZIsZvL+SpI5DSiAByDX6B4V4YdLz81XZ1l6fSQT6WL1ACc41Dq/xT71fpMfZ/VCPOJ5HZOHy+H
G+TdQWBHyjb/Xs8dMZc8k+xw2CBaxy9DLY/CRxTMl86FO5ZpAl06toXjmG+fhoBwlJnJhIQRWAKm
V1dVeVcLTYyNotDpQOb7iSzvRCb5holoRi1pUq5+R4OjBclBAGg2/oxZiGeN/D8yGNR1c2mSRLcn
5g+kTGtzWQ/Jx/a5Qm1jPb+ELDLdPsBr+hivWVfPy6IMPBOfsK790pJh6aa9NCUv8BFegDrCAiQ9
EOfE8qp9VKZdzjBC01710xKE4piU5NxGA5cRGKg+DKbhHDDoLBdXv7oj0yg81+TIFnpddd1wiJYw
TBPiXa+gXZtMKKPwCTd73j9IJf5xYPDRobNKpvMsGvBzuKpE9reSubSrYVROuN0le6dE0pmCy12I
honkXijh7j18AAiVAszixrpazsccSjwM+KvIYp/hWZTqSxG5EavbO8MFR40tlTVc7zT2wLt2bBQJ
ZPwY0TTY/MG56ao+iGRQcCjnNXbfERm7EHmJ7vMzW13ThSduyJm0ZHbvS3yHEe5IFH09qmt2Spyf
GkB0U367yfRVmzVIujsD3AwWCe0/qyTEpTd688eMwgGRK1h8d3yLDMLB6ERO7L0aHiEBcKrIHCzO
bdn0o3pP/Lxjo8DjcHlhGGusaHNQjqrwryGcZwRc9ipU1p4YaULStEB5pTFSmH5UJQIyDnx9Xyy2
jlmyn9SNzKb1rBBhGCOzJtmmvxYbKnExmtqbyQbvu4ZSogToAXGjlLlFOGLFaaLBI54Y7PbyDffV
zLT2pA1qnU3KUSrZKwz9U2MEPc5pgNLbeR5UutTs4ldTQ7SiqBVy8+RKKQE8VND11ZkgHdg/AfXH
cFH4NJ1UZ/MBG4n0Mrzs3oHsYheBcp0mnR8jXTNrOKYmYm4A3EHkNI/DjAKRMuPe+Eq4ztNTGCX0
fhGusapVRmYdU4k4t/v5c0uUr39kCZ/98SXMV5wSWpM/gPn9SG2EYAYSckdZCYfOUUCcotUpeOzO
3i3nvvetFa74M5Jda3YXzLz80bNOMm5Gqb547RmyGsIH43MpewgWT7d2emN8+JrsX9QNKcg/4RI1
sKTBJGLbexW7MSM/MhbLxuwqU559WBgJ7dl2dYJIhJK57cjAKlVB5KKrSsJuccEfgrmejfZoxtN7
wfxzQ6wQK0FjclG8M6yBASqSR3apPFi7nC6PEbRjwIq6+e0SwtaYXORbjuDkPP6+iT82UC7gbucl
CgvB3z9cwzB1XmMqkTXM4ei+/Uky70AMT0PMGsuodfUwqaUACbf4OpwEXDXUAiws//v/cnGnxKFs
s9Y0cbU15O7yPTmLxFDgCCPKRO6ICyj0Ji+xTxTNvLtBcxuqSfPkhsrjS+eSCycBn8IE6mUAQpWK
HqMcjTNx+tMP/i2EWYa/EvClopPmSSSfk7PrZu1Cfm+Q4mbrSQHsBVXVGrCIqzw45N9MYBeFD/4U
2POWyERtHOaGEY/CISK38F39x28aYc+DmiWVGdmvZ7yVzxhPV5ZoQ5YQ2kFU0V7hJ91XUYzbkg0V
9GTh5Pes/bSTHyH23WAlfXAW+a9lKu+QbVTFqsgz0BG68XD37H+AgDVfS76MwF/Faz7P511XCLA5
tFgQLY4CJyQKNcnhD2VkHwT7WykPxvLEaPPb0m+oQYHCtJ0VHt9T6l6VRAoGMc6O8LZETKNIR5dF
0Nh0PsUkKjZ6DElJvHbvIe69QQ39DouIEhPtrzYgAu/jkiRyWDmTfuF6TwCDsEyz6v/0ovBTtgDe
6SG6MGM0raPW7nnN7JD2VTEoa7k5xSuAk9dTuB0bGCheMEmmbfsIZDvI9FBG30qO9iAG7CUdikht
bK8PKGSOb/6pbPtWbThiAS/DvJT5dOSf/9+M8qy7PSIAB7DlfeAB+4w+i+tEIpy+LAB3D8H8kI5K
rVOnMJjfEV4TmZ2pmsrqaVou3ORSMV50TpJ3U1LTllm0hdtkhcmWKbHKnyYZGr5hd+/rbKtTCMK+
cMsKf9jXi5AVbBAlBYl+3Ec3OOd1vheEr7qsas3DvXmdaof/L29pqZdcRg+G+o3p8mNIlTfX1gql
ieTEB9zTw8DrwDnT2S/YnpX2svHmGVtHNU8SKHwkxP1fUeerbmBX4OrSsoESGF5ZAisEpHtnF9nI
Mf4Uf2zTxQAFV044sjtC8ukwnIX6ttVwMKq5b3MI9UBdjyDSNNEsYUEo/UsMtHJtv7RdIYWzK3NW
3uXWcIdc+sWfMPaFgxh77wYJj13hJJIDUPTI8eFOyM8pvHnI2d5++FXpGYMstVKiPrw6Bml5qkmT
sLVIj0+CCb7dV1vnEfwdCzQMUsELwYYfr5kLYD1NIivVyQFhuOFQb3BcW4bF/EXUsWIylN4702MV
+ld8MP3jUw6nrlsbV81484ilMgqSsBoIqOHCWpaHqkls4wj1ijs0jvkUFQJEsFzrrzCTZHZB9Ahf
101RhYQ19L+RxnuDrBzKn1QQ4/RA0sTOGfC5sRllmlRUypyBG+nssGxWNtsndqLB/8ga+XY3xjKH
wdWNf29YKhJ07bUJN1WUq3JFMzw1th49RvQsjXYHMmfBVYKQ4aO6MA70u2c+NHqsUlZfAabKEPKn
BgnXAAW4h+tLZEJYjLlrYmcfPc3VOkSMfSE1OAwiVVtVCeumCGcar1E31TdKYIfEkr8n/pwtj7JM
CULMnrOimgscmHJbevSGVfWaw1fTanyq+5HEW063+JmhA2pT70uXMIZY4oB2Ox+DdW/7sUNSICYR
Nht5mwk0aaTAat35Yq9aA5VyVVNo8GynnRmZ1VlAkS9Orkdbs1WE6zxciXlMHR2dh8H/Qi2qDHQa
TlyM4Sbs813ZBe448ZPfnTo7uYj8rHq3awkAXg5LnMkOCaBYXaTtXTPVDYwGx9quV3CKYvO56KX8
lj3Fg+JjTlI6UsgKhtCFTPtDG4vJAdzwEHB5e/2ofl0ZI+F3SgsgNQLzXjw+LfmIzyYCMFxqF4EU
1C3+TV2sQVN3vBn/r273CBpDVK9yQ8WcvHlmwzckSeyphbwXuSW9XKVi6nCWXowdtpfP9vqv/Ven
ef05C0NPI0DDP/cuklcKcl9f+2WEsznUcwMilEgh58jYFHahb6G4WMsafHde3zZbqOXVS7mVnlSv
idJzJef1sw0YlXKaUzdVIxNqa8RRV4DwxhhXGhgWNYsvRUuLGmJdS9wZjZJ/+qdgMQdxXxQllY4S
78T7CpygcQxWpZ9SivQr/LZsVUyj5WRdeUIgprwbFmm5OI8q+E6C24o+iZnKMQNKnIMsV6IdYhr5
bDvIqT/bTbmo1hL2k5O2jMb0Ucx64pXlusgdv3BxLFuNRbRpwiMi1hiuOOlLC8xfXXIt9Q0JKz6I
hbKD51JgCTO2LB0b3qVdItaS+R+JH+Nkm+w6DeWD7l8xIg4sh7jmUt7DxQzgtTqNoCNLPqR4khY6
eHGEmOdG/zGUuf9dEXhEiLdgPMNsmw6+A7HmQ4gf/RZV5j7Dqf7lh9ydCPtyri6UsUBv1D81TXAf
QYboIrMuiap1K8DGbtwhFfF2lt+94QlTyImFCmevGVUcE31awCkuiG703Ofc+E+zwTu6Q5aJlkby
yTf1ph04s2D4Ht0hFnbi8j92w3HjUFdrx2O89Dph4nV1EzULKiRB8Z1geNcLPDFpTZpK0IH7FFHb
/BF4x4OMNJikbbUHDVQYTDZFzJTNp17sCR5AXmMZ10EvhrL4TWiRu0fqPOtvC1YaJF4AO8aBpX0r
v78MfY2+FzCZx8jQd6JKWxknIZkoGj4fdIgLaSzrkBEZBujrABm3I/hhsB8ZB/v7UIdxpOt6B/Eh
D1Fg80z2ThqumFV73+zc2By1l1OYXR8avCZW3KJFEcs4fOVHhGQpGKpZzEQLbnZ6CdxzS8WTrJTn
F7rbpjRhAu5kjSQhUHU2RQBsz1nMZ39eYRxo8ZUzBWVPWO8hnYPbM9Oq4wbjJzzV3CkcJNafG5us
9GAAgT5Ec2QnWQKefIiuKq84ehXQehcOj7TUItrnu0yDmFn6tNyzRAzfeL/s3H+lS42XCSenggd9
wyiqIb6tDATOGjafY/hiQ+kK4abdxM0qb2XhmxUFaOzb07XZDxv3iK5kMmT0hoRpek0TSm88Mbgv
2B9nawEQjLj0SW94FziQZzMtMnGOqq+VWe/fByhNmN41qmnlVvzjMhvvGkrQhJhz0+x30WFaxNKC
SM2fFmjzYT6QGSk3ElAaB+irAKVO9KJpz0/Ylc3KUiAV2Yq0Y1U2N2hv0NVtqn7Ce0MWoHpMaVyK
T39+bvyaXBSBN29nONb+v97TPHz0PKTME+wrz4iWbfhZ1crOh7FAt4ZAUsf05xcBnsynf8NaOO00
EloUjvb7pxXtC9uKeOrVfekUoVZHYh9W3erFPpJsvuBSRnQ1RFFuyk7zy0zQyaS7ZAmrKdaD1N4C
bkGIVQJRhaZ/zmJwZRZFb8/Da4tK9tg2T58Qap2eRyFUHksPVj0VC65aoJn7WSyqb2IGXe8InGwt
R3Z3udEUHsBP987zw5znlBNk37fThM6mBFssMPxc9cxw4TM86FGrlAYFfdhsiNWH59OMSF2QY8U7
83G8Q5SbMxZ0V8aYrn8CeCEr/kO+N1af0M4AmvqLoY/m1a+xmy5Enz1QQmKYSjKuQ7tlWvLxeF6a
/RYnA1Sq60QowiLVoZDi56ySnWmgs392Rfvu+PCJejD79rGGPMopvILShz7jaowuPD5exlthIFRw
2wd1ZwFYxJXCUZmS8eFNMrfP5LVlXbeuzLBnfHclfPstWpsJyKDW6BBLS73RvKWYCzhVXZqkmXzU
4nqwESHwuQ+Muz+Spo6yOyNLmgm5RTKlj9M7QSPikDECDlP1n/3hHZmtXH7bJEtjknUQtimFbICT
xULFKG6llX9bwIQMk14CmuVnYcY+I2HveFD7mVNywiVvv+TrSpYLiGUd+BJu+CfHPUhhgYsRwq6O
kd5aVjmhQEO7Bm8Z+muvfcxjie1kj39J3VkRtUeKMqqVYjEh2c9QLZWKsNPthgLRWmrGMkESPgAK
xtw7KJDFUtkmHqOKqZyhAW9mXwG8gU5WrUKTh2a7L1E9regfqy83uuZ1r5WErTFZ43ymHDulr9Q9
+QYQYAFf8zU833pzcJ1DL3bl3sUan79D0PqcuXSJAXohVpKESrVORruQgznTKFR4a/w1aYBWG9J7
HfDxFbsmnGCi3GOqMJVJzO/Bg14AwyJ4l5NCRXPw4+JeuF4J7rIcUXZFvLMXzDI9k14T0wsdEAJM
SodBbwn07ES/CwV6KPH2fh0GEWbolx2rX/LRPc/Dx3FcLpbLKw2x5KxnQCQ93QvnGbQy09VcQ6XV
LQwvwDiRsHmH9jJ7SzXLMfVKZL313YDE0YE2/OixJ7wHjxJi1GyBXdyQv9hL0KRGZkFHDvttXx8v
vkp4Yi5QCUHaqAlIsRrw1FkEyh27BkFSHe8vGO5Qvr0HdXABJ73nBI0X1C+30i6ABkiBjuK84aSL
kV70XF7cYQqUXua8HYk+kxbBikO29Rb5gmmBh4nq9BaZOP81KJJRL2vTt52EJlMhjkm3Eh0L81TS
YIaiVcr4tSyFaPAm1jmSy60O6nG0VjpP72rDYdg1R/kDiW4YAuBt+3Zq+ZQ4elSY6XCH0K972JSD
jLIjz3k3SS59gB2+gm/BGu+xdkE1auTTh9fYezGqmATyId64L0g+z6cTGQmpmuUetZn28swLaev1
stGDtGj/2PZleJajuszP/MivsrOnkY+Fy7O/tzQQZK4Klr4IUN8cYI9bycrig4RYLUwUXZcODQNx
UzKNBcVXzxDWoMZMAZFG9doy799dq8l15Na3PpyPKoV9qglK1K5gYPAXDiPKF3EeU/+8jCKqdI9w
LI6fkKswjSGDG3UzTyA1/8oj6pdLlc2zwkEzHQBbMDLuzYbXsAuIUKCgrmiS+tscnywHhyc/npIJ
b3dXHF8ble05qnlsha1i7SNUqECkd/EFBLVc8IkBbRR6Xb7Vy/J1eMh+lgL/4jbITJMzMFGQ7pSR
uqjA3f2MkHaehKuYZ+iu9XdQgdWBu1Lf5VPKSXe5SD+g3pYQhq1TRLMoMfnKt2Wg1wIQyE68RGQE
uDdKCNaitfriP7OJew6zB4X+jYMenbEZu9x+Pvin7QHozINmj54o+udRqPg/DInWwctZ9Vbqrtbo
rb/Xavmc72rKv/xRhhOAx6G2Pe8mvzz/oP9GeEyPmyaoeeA7qnNPly1sex/04XN48sZ/Vj9UZxMc
X2Znk0M87+tVouWy86tqxvmb8rztD/lFY58QPGXAfN9cchRXBf4Wy8T1z501LnXwHpLp4p9Ko9ZC
e3H3rQUKbwm5+tX9/04BnbM59t4ZPba6cX1B8PEA7CGcw5SGB7XaA1kU5VX5gYzKg/Npju2xiNKr
wHtBdpmX7A91llbPQogVS2jLFpMkp9+RNqOQZzDSRIpgtIwD3RrJcSwFBuOW6Uz7VMEkrbdnF+26
bbBKsc1bVI4VMTozemueLky+cgaWr4M3cMtXhsiM3Y7fzdwoKgqsXOMgxN8DjUrU+1rNdK90xYja
cA5bGuH+XgjL1xXjA53EtMNjN60zkik1m3OaBHWCU7lI5mVIl5Abt9PYkkhrRQekVfVJYXnzv9LL
2nl2jvRF7GJJxZUjA6TI9AKxtGKxXI6zT7cbfgymZci9z94caDxkatldbUeXLTDeluEN8hgczh80
RFKnagtBFmjxL0FS39enUEZAEjImTOlxk1PwdVWATm6IaBdsHE/nPKLz0h0A20WUKxJWENL/8CsH
3TmqnHjLyFWvdW9YfMvN8Bxl/XzNfBUAG37QCILt7IzbalWih0DGs5b4AdgGYnGh7jFvGL0FQ9J3
uj25Eq8Uq64jXJHmMoiiNKcqodWiTvGB0GhpYZuzYsq/gB7gPT6z4MULcChzkhjFbPToYdy/ct0C
w6Xv0RyHqlmUdntigMYI9ILtXt6UpGH+ieu27YaH00HprXKsSzemFEAkeBGMOHML/K5uyJ0PPWWN
VgTifghaugPVDkgvpEy7okQay4e2hzlTJzIipHTB6WL/ANnPWeoAkq2vTCTOkBv8Qt0wl0QVchmN
EnZJkfavnhGII9JrP4pqSJXpuWO40ZUqfhBzkMakos88Aacd8ZIqginYc5vf/FH1j6OB3/joiQkh
YZGbK7d1rZ72TfbI7CeC1LT3nmfSRs6YGNxcpSn5aicwIjG2CM7+9RXavD4bkswKOkmDnXpFHpDa
AImLyR8qH9/tmOYQwKEHYVXWi23CW2agaz8awnca7DaMvSgpalf83cMiLIX2+p7FjHEDacoQzO4x
p6jP6Yj92Flg72pF2dHlikAOfVE9KIvvsVuyWOqwd4f5XcS9D9R6APGdYFIY6Dmry8zPIrhuXJfC
6q/LSdQO4vtEMu7csbN88rAku1B9hmEscQMf2IIz9VJ4MUJYX8n6VaAl+H90kF+EuHjfHss1P2va
0w13U59iMtS3mLgO3/rYkfJjIgF7dCWoJRa10Y/sThugnUDTMORJw5zm+gPo2rtMi4jlbjnqlAQU
8UWoK3/fiTfkA+5PY/vzGeXtHy/jj9kSXGmcbvyGcYlKp6zNk1ALaxR2Y9VZgMFeBp/X3um3d8mA
1SvN00u3xcSfU3HsjKeRheKcfd5WTuN5EPXsXbGSxlYHgEQMA91htmPjdi1888+7ZOGx4duhfbU+
2Y39Fku+gzexkmL4ySNdvWDkdi0o/HaMIzOHly8OknmkiA+LV2uKNlvP0dEsarESR7gyMvoRZgxk
YymqQo2kxnvEA5Axnl0yA12SeKt4esUt5pdtSpthZTxWumOyAJSVhHq8JHCxRUz+om2TH97ZNR/3
90rwxyD0LhQm+sNy6n0XQmQAwUnndRuQtmdvuozFqvcH5tIp/ye+piiVdSqJMOqKl3jDlgkWgUxV
OSa5IKGisY7rDGD+zERrMBlxcKOItwE00XoOY7pGmhCHsyTKEwnuCAXNrMc25Np3btNIneAo4VLD
2q9ku+nOs1bO8ObHJqsTNUMSA+XAoyAYHbNy0jG8qqNgLaDF+q3cYjHhJJn9WAobDW/fGtdVBIk5
LQyWT/AAxqeTRjusXhd9t7m55Wx06xevhKalj4gBsXm5WpbInlEDrFJKFaR5a9WhFlaUelRpa8Ea
O/AGwpMDZHKvcYBe+byn2lALVGLebD+rEX9UNEHUqKcyj+fJpY0CeXnDUBzXKuQj2kZV6br4YwFs
CpRs8UUlxApNlL/wnTqNmaqy28OHQ2jlGZ+TzY6pqyCoV4XvRaD1b7XipmcqoCyahot2cXRPw5jM
VIeBQ27TL52TInNO1ix/ahRRfDohPvMRljgdbzplweGJfSuyiz2/+l2DN37QNGhdf5kA+Hr7kNex
aeEx0cMUBiPEfFn/0hJArxzuGhBI88wW2a1KDFHbdrwtyML4iKcsNiM+DW6mSbpSfEOtUlD15+aL
7def+8EsxK2npXnwg3uGtELyJCtnA1qWs8M4b/bGbTmAuL7yLai/T8uC/TknXgr7TqS6hZUom8No
8WlSQbHuKwtdiH5RSjIixb5Glx5JKygqQYnrwGzQ7klbbeoFCktgDMdD63pLiS0M/mh99TqA1k83
DFQ17sLRKDjTWZFDPV797aKDYQHpHxRh9B1i7HNUgalULw+lyyPmwhYjILJZGRnNy2yJePimikFw
hu/qUs3eZ0IX464VCDe8Ptv9Ih3ibMJEDEgR+bl3Bv5K5+AiEVEeC+MT6FjmDU2nWHCYvCL97FiP
Id5V3Gt8eFa34DKtf2Nvl0YaEbVd6zTVb5+RneIeNb3MiVFah7Kf7X4IM62GUkFTwQEl/1wNc344
KJxewXFHrk+PLC32R7xOQg/flJdcenQ2reQK1arKcHYSni2f4OZHfUplyi3DtMV7OolIG/87CLDB
Gzmol0kDhdqtAuhGz81r3TmzKW69fPUDciih3sUVio6+nzkYdV7aZlRGu5Ak5fWrV9EgbM/9jVZ0
hT4t9HXoRN5Vu28IMcobxRqDMFNYCqGFt+pEbuX3KF7HFGv82tzWQMb/12g+DOtAZEKSxsYvKYf1
RNni4wDrMx1s3yK9BckJLvIKD/9iWCq8BlmVlVN99MkqdLQcV7WcMLTtFtboJmNnbeRXL59Q4iCa
7wqgIJWNzgnSS4wn2KWzg3gEAUaTU/W/2Hy3XIey3jHC+YgwJD6dSUPO2p5uF5HZWFMSqZKX9Mpl
2WGYJt6w/XmhBvCOvznr8ztuy4kdV835gueGL27UWlp8qsCo7TGnmi1KVchfQyTKsfsazkWek31Z
7Rl1lflUfHntubz+VY2oRC/2446r29KumhlU3NEaeHQCgMFPuiTQ60SHphaHNrSng1pK4Rl3HvuL
KX0mRaC3Gky7LEfjcQ+BHdheATdOSsATnKZrBW1wNk1M94X/tFvdK/9tSkVqI5/x+FkD7HTE5826
ur1z1zT5IEVXdwGKRGXg0L4WKpHKan7csJCcUx5CMru7Yv7b8LPfig4QS4rwdE50TrWuxq7boKJg
Y2kYyj/SKaDEERyGN7MYdZVP9tLzrHUbCWYmwA3OH8TNAcqjldCmDH9zbUqZl5KPrhvXE0X+4PIw
CMxwSJiCC5qMbx33CmOT1x4SVGKQjnMa84Hy4fjy90F/5jWTeN/FqhpnrOJ+jA9TeYp3mTUb+AtM
1rKRtqBKFAtGq4uCKDob3fS6Qad9ye8RNwNbgt70KOgA6cEmKMGiqJsZRvWTaA1DHLg6+MHB+3NM
COoD1NDTeOpmTtEI8DOuYV1iBRbSlUvLzz/7VyvA0Pt+u3DENINxnoYvFkK8vHoW+//YOONrwn3x
QAupG9LQAfwEJ7HmEcOL5cqzKFRHNwHgfXEUrfkosbK+rOWmMi2vI6cumf6ejowabn9np8Cj68/W
eQ/ukmPzdi27ng23fHWcln4AhqtbuEX7fffWQR4+VyR87LEfq6+h0XKdpKOc2vJMdZC+wHK9zPGr
QRud1yb45zbKQIGue06doo2thXV6sCHogctvsrU78YfqyLaHdhPz77HbMBgaGAxdKKlu6XLr89G8
asxsnboqV7pUb81zIzJAUl/tAKT1ZPQl9ic9Ga0OzhvUzsGNGs3E3ShCvEArcC6FqJ1957ptLieP
5WALWIf4YWWFKHNJ6lb6/Cmu5kBinWZ3So8SNJ7AZkPp87L7AoBwmtJ0F//58734Y51MEE/vVIsZ
vheNMb+NqCmJ4z7ephYyROC82oY6tSTD35MGzB4UcQOUjym4xgY/S39QNhvQcEnRm3VocEWhIv9X
BtM2Wja9Sy9wfWmKyf3Aomts+jRA5jh56zdpB8MCMr117H56S+r0R4LKOtucezqKKuXiHfXysOFd
r2ZUWAgzCmYtdjB1fmX4ZLudKIWMlThjwszD8IHy0lPHz9NkButipkAZFvLmg21M7oUpthvhTpYL
42WWYlfZ/RhOP4XwofWeV7P4LNwDJNSj/U+RBVMZi/Np0Qzcq6eOtPWZJbBo1B6tvVL1To3k2Rvl
lbJKOFeSZS6jxL2JLezNhQy6nwzewJk/1uTlIIeqvdpfWZgW6BEY/zQ/RRIkKFABjrH7ZR77xWJs
3w+Xpu3mE0/FKctxuS2rz1SRdVNXOjLQeRJstRu0rMlLTVp06w2TZDRNrXkkmG31x2nojwkBCl2i
QtYt6zGwWquhEyaEMu4GfScYCM7UhvnhSR1V3RirlyfbuskJd6n8MKSzXdNalO347poTHfzpK5yZ
YsA1xlOyQuE9QiK5+M9sOfleWoKDs5RL6htk1+QHDLUuovGwyos9ZLOrza1ilBWNXlusQNnUQBi1
VLSK5jWX5ik0Q1pk3/fZcJoTsh/UDHbzv3g7+C7M45FtB0UTtT57/nFnC4VLxH23vbGeg6M+BoXO
pX2p9WmtPmL2RBiwevzzL0rsEhdUTGZyVNUoXIf8qQJPTkHSf6Cp6vFboTzwjooxnAiSnE2IfjyI
PUyTBLfnIauji0/NqtOb0MG1329J57AI/EtHFCcdQafGz7bALAAbikZtx2rV2n1Xi4hG9fMbrscM
z9SMR6C54Cj6051y+xo3ha+ZlEoT7CTB0ChyusYmGrz5/AlfE6kV6k/Ske0UqhItQ6vXby4LUvaA
eBWIAmV3yn6Mq/ZyxIfukw1o7EvD7JbiZykpIqWvJgQt4JTQFvN9adzylQK9TpcRZHxe8/LRtRAe
HMKK+VifUKP2m2yEKMipZ5F5Jsw9jHAndl7E+GsiO5x5nY4SSN8z1c0rNeTXFDiBvxXQdpAYVMd3
vR9IEBPI2dGftPkwoc5jfhPlgw68Pe8169hKOVdGzLE3IGwVjZR7NPldkUMhGsbxKPB0tOuji47e
we5VcYnJm/0vMCh7hpDijBuC4QcWzNYw3hjURy/KCileCcavIwmzvzG2j8yJRe8yeIQcoqV7oBfA
fpqcXUY61HMzVi+C3jOaaPIY4NTp7XN2pye9EBxDtd0g0IieI4iy0E7ivP+5i41km4/tVqHCHkjD
5TpFtwqiShe8AGahDf/LhnbdPSpXcinV2OxhSIpn0vXKRDsW4P/Nj3YVmOdEbyUGldp+CapqwCgJ
c6lCl8bLAaFOD2+kgQf7GuxLswga8QJXM3Njs+J37H3WhJI/pxSP6Oe6yP9endjDc7G478iUfUKC
owwpS9TkU2VDFi/wG11TyIXd0l+aQkd2JXng2lQ76XoMqNDUoSSNjuCI9uL36QQWn5BNPznbS96b
rKdUcTn4NqcQGeRgEBReLAKSVtxZgPkoPfLUngN/7c3/g8Y2B72/wX/jKqskxTt5/wUK252yil9L
UTVGhV1eiGc6bgrL6vksLAhEGkDa58uO20KgBEXOWalCJ0El/MvB6/x0o7e9hwLv+MT4tDIMxh8W
U/Rxd2N3/qWmgzPS5OQ/7O9KLs5SZUy/jjAJPch2TB+Z/LBdaA56UelEdB+zCV6XXU9VMUe2NRIL
3LEaDJ+WKdssSpFMME7btBruPE/vSWImnx8ChHnTwq6wnroklhcpFLbF8pA6U/J/yX/ctp2RIXFi
isRTjGbUnBicTyWbz+qQrYYbhBjnvNNVHgYrPRpWTN7/QiMgj1nxoqQqrB/W+FZDnoW50/m9ZjXC
ZJ3uHfDR0jAKRc/Ao5q4l6Wyt+WscN+/axzs5ZorrDiQnJz6fAYSptMLBmUnCCW56n8e/jOdOvUG
cZQIpjCNNjGn261G3GXVY/0TjPjsSINl0+JixF6MJi694T8XFFUSNwNmmrVJd7UlE0osJ6yhqOLU
Er6xVk+jY64HKw13IxPDTNGQ8U/imgHkEmAaaw4jS5JSqKrkYIwLh7ecgeRFa/5IGVyMvfr7HGMG
uSGpRcRy03TpLpnSQnuFdannwlJLw12hf9JcQN0BDL9PdmiohvQLea1bxgU6kPQWHsclt7uZqzRQ
JZL6ZHyTtkwI3qGLYyWFzz87H8ZTzHk2JyaAfbmYpSZLveF5LAWSTZU9f63HVbczvrhcFF/mg+PW
arO2gqEi4IpykYWROmmQm96qKtFKvEwKdUwbf9hKANSqNF2QZuVrLZBsrI/+IEWFdlN5PSIg8aGp
/v4u08LxqwyzciE0z9Am/nWUn5CJ/I2zIJhhufi73pn1Nw3z8CEn9oxBtKZ4N5Q6RBgV4PROTehs
rv43E0hWCx5NxJVvPGpGAyZKqCqtDLU+didu0cAb5rDlt9W2cfQQ+r15C0009SD75L914KMMBKwI
7t8kMqzF6ZiVcuRCQXOiHRr2uWlMAVuUJyl1ECV6EYiYbZOB5OmRkQ1OCFPwgX3XWe+fxReX6r6R
x/AslVzKVU0KV/xovPF0E5X3ozS/B3etksdG0jTE40g01tPApwrY/4kFm90RjUVbygAg0++gjVl1
KrrJ3n8qN2B6twKYrBX9otA3ye1R0798j14hCUPgPhtwNj0zxQnyjBOCkWG2o6Xf2NXFAjqBsNSz
hvLUFAx9VPoEsKOvIWSzfNuKPmok84HfMnrpVaCVKHAljmZtWOV4Yqh40tmxmmQ6SKdN1/0Bvsbw
+WuQbk4sRKFXphfKifha7mha4KZCxm0KTqrf3aekNoex1/xBwu3UZkjhpWqutV9Kg+se+upNEMYx
mPp6JVNe0zCCe6jFlJnM4a98xNlrql2kWugTyPfPynZzD+zw4oTnLCBxq9RtsDMArv57KD3pjhb+
tKe+DKXPcXPyu+8sm+bbyma/xLL60xggiZs2HFFC9xV4AfFRKT5QhgJfElQjDZJ/o2IerRQXE07l
RBqJLVNP+0lSWbWlTXVCBJZup1DpfDo5/7eoJYCrVE49uA110IPoIihb7qda1qeGK96uRJ7FcUDe
Q7/dOPf/UMLchESt5rC4MdrHX/uwz7D2srwmHDmDDZoQ3Lv7UN7VOPTEUoXBRhgGo6HU65fw/w/K
Ormy4OQcYud0b82+IuHuppOsGraslDLNldrZBf8tz3CkVteQzOzPcgcqCi/GgSvbCFrkzJlRl2ws
Bqu0hXR52MBFjgVtl9aQyfCkZLfSoWtYVL/0qBbyfJiEEMmdl9y1UDKB+8RHYwJngqS19Xj0oBOh
K8VHAuk90w8oAfNcmAVSsGran+4g0lp21Glglx3JvT+ohgzs1EwIxkeo1yKbFrhT7RDhhEtmrhsH
EV1uCZov8wlhJ3E+HuDe2lBPxSaYRMITsPnDfbIvKmEwaVPXQRluEqhxlNHDED1EvxSgirAlYJ/o
3C6S8/CMHBdDvn0WvEO+z4deKnhXVFTWNcjBzOWQ8ypg5vZSQ+AsPlkGrVWOs2dUedFI19M5czSd
3XrUP/n4pV/GmV8lUAoVYxknfhCHpogB4Pc+54frthmtee1rsbsZqz5Pp5SL9IzmXcvKEG4CgBbs
y4d9jtjc9MxyYSAC6N8E7S4mNBbLazH4y2du4XDbdwp+1ULr6KPpZz7J+xjawthCVEwtWJkg2b0a
AUZwniOw1gkKMy6RNfKwPDte3UvEZ+82wSf/urRbGtWkTYH49nABa8PphPyYd9SRlSQTtHo3PM4f
0wj8MhsHRNQGxxddADtmpafPPKXdXLvu5be3Vewwm7NMJ+ueRef5vpiF8jKxtRn7IKQ8kRg0ctiC
CUwYzp+oY4c0ahXUFxPjA1LIYbDY7SUz2IdliaPrlsjfbPCO0JkRgS8DSOmVHmhCJ3PabaCMQGYJ
8kimga/ler7iiuGVH6kCJpJLaoFsKuNng17uNNmB631r1uat28LeXzopuOvKPa/rzuBwYodnsRD+
lZz3yCXKbnL4WNpJ88H3r87ztfGjbHNiFlTxsVVxVykYWNMyyrZnUl6ARlc1yvzr0HCEt+3L0foj
70cIQCKk6SubNVwJjst//fYlfwJYvqDFeGNgB2V6t+edvy4aAynovD1+lZmeGk3GfvXfUXBJ43O8
wwKOOq7Taxd3iKZ+B5+GP1UhbMhFHYDSA3TKhOKLw/RdKdNZwDxY3cdRN46m2ZklcbVTrffLHDkz
IIEeIJZfue+SHHCsyL9AlVR2CAt2L5UP4aOT+uBKoKDgvr4sZ4TEgUFx9LMOxQzmBHsSzCWkVEq4
nMMLVDxpr4So5n1+P/YZJFc8c+Osj+0VBjz22MwaPlrkrQmxXD2wA+mftTXcH1st1HrO9Q4+rY+V
xKGQtrKgt2MaEKnQDQ4QiN4rDEiOOCoLfGJGFLMrCOVXV6xNUF9SePPuD18yp9VIDZ4qzy34vslM
zKiZOHXFV8ER/HtBkaA06Hu02gHROqdh7SJ3R0fwD1i2BJZyA1XzW626hfxK/zWoafc2lTp4cv+o
0gFwSeTGs1+eGdXel1I1cz1iO8zOWSzXFN32nFhxIvIIWtliDS9P/dNBtXLWtAdWoovE5d+0w7nU
FWAcY8UFUXUc0s+6ARhroTiBx6PkVGHzhqcl8lafNuNrdvYFEIqe0/K0b7uOPwL+L6X4ApNby6OG
6+Mn2nn+Kra61z56GfKYaEMWSA1MjHLIBecIYCMZVLUwQ2HgKWyZgToq0q7s10F90pIo2MaHIiOZ
NbHXCcWRSHts2l3E42sYtrSjn3H2g5TTa0/hFCMMZs7MBxbNFXE9FPqBPcorqzcVObGz9DKZ+ldM
yEvFOdpjPuIq3FwhHtOtVLt4ddmdamUFwI37JqV6y6XMPizR0fsutSl9n7DaXIsMNeY44BP8XI5j
WbBqGKJ2GrFiWEHR5DxvFJbEbNdw7k9fnDuuESRZujrhkwlhAQWePxDeJjorMqMAdIdYVRUDPZ6G
0pEQ2y+OnYMfjNXEAue4tVbQIJWIU7v6IaMwK4pYje+sMHl5dNqREbXw1+6qeKJQ91xREJLP+6LW
GMDCUq/h/rNikF1RwenCOQ0dCTaoFF2BfKv4JENKW/y+aD7PiZOX2yf24apcl/9B/fk+DLWylWui
ccsIYptDBDIA38dfcpjG3lA/36EO3WrvixYIdygPq6WjPHffQkyoh/+AAt+6v8zxvKvpr7kV8IbW
wNIdWXqoUfUbSuQkNnY/t39pW7O7RPA7qFfEa/+KYhTnunXeTGyK/b4YZIup+ZgplhZVYOzb25G0
xYygPWZ10IwWZmOWPfasbKka8JTy8erUje8bfoj7MDnKG9nhDwC16qBCHrEjRsnI85Ca4MtqQT1V
vLGJBhbnA/SkIv3f+J8EGFIOtx4fT9ywqV+j6UASmn0tCIjxe3lxszyaYopmy5s/o1m8j39VnWbz
H5SeTouoxUNW2DZE85B4wijBHW3ZwM4Ptd51fa6ktVOpKup4+YRbouOKOKJTRaOX2QpUq8Eu59Ce
qaFZ6P8Qa1oRkZ6OVP/D4f1D0jDV0lwHkzPb4yexVHdstjwG0tdFH+WYqsWI9c56iA7ZgsiRaF14
P4mGiKIW4WFpByAKXOgMc1l2hgTdwVdWN0YIlJ9OledTYdCxWhPOLryWcu/aLBm313nNmO8V73oH
2sbH8lOe+zIrUHPvzwK9lMFZt9QWLPhdrbmrIV44kUvjxu1RuLssCvX2RqOkYKLtisCtI62r7wIG
cPsRD76XPHdn37GRgLvkfYTVnSvezL2FfHRh3bg1gcU/ExN0DMQoo/kcYx7y5y4vUe3LAdyZ43IV
w4KYlQBn8McmJSxU7gHcZe6CtL4IuZf0OFVcWDiiVyMXhIn+VrdoB8dTbLE+1lZ9DMqsJV1CNYiX
BlZgdwWagA1hL2xhJDAZRyfpTuHOp2zns5ZUDYPIL3UW/05/uI9+kSm3fUbucfDRbCha1css4Hc3
Tw1DeHa2C90N5z5QT0kniTY2W2e/9wjih7IqptKvUfZx39yKhcbamxu9rgdyTsoT1xzZ2lrAEjXP
e7WFxTgrBjIKfs/waMQX7ljqRU05MuQYAVaUpGw3mBO7O4ttIvJFJXtX6+t6Mn40RuRqnJ0B86d/
Kdi6ippr8HTIXhZz6npN3l5Q/Lxi623Te7wQtLbLnQyiivSl7XOs0bKIoHNKoualbISOAYfWmbqi
kws/urlSq/KCDAkf3gZgDejFOgsxhsqaH0UCHIhmimJDsyHNpClFRIU8Rv3EXlJDi+/kJ8bZx+T8
k3veOgzxwswG8246OfHCOiFJK5NTHgekcRt/g1EJD3FSYl0Fib8OlQL9D7zj2Y29u+cyNVG4a1pj
swchOV1W0ADd1ZtO2UaBTdFXp26msOIJH9i7FR+t4ht6MViVJ5mAoyTYm/xxNHFKDjF2VFC+jGd+
6kWOqBOQKdSJt0X4dJC0PDkUM6r4K55zJvLstSJzrR91ku+bXIPXxLU1X3ceHoIKDTOXz0ZdCM9j
Av2L1pj0I9OX6971RjoRtg/OHS3Wz+tjX4jnQY1RU7XLHNGODPxBeFJDMvbrlvGf/qLuljFH3gsz
6eFI6sxOf1gjYa0MFWsu+YpCEyHicsCMrMklpYWmH6vCDA5t4CbkCtovuw/C1D9GU3vKbmK1sFKq
hb2qejdtv7hEwJEU6mN6v60pr70YJdC3Ty1JAnvOKeIpez4Ax2rATcP8IpASyOLNU16FbLJVFjZd
Fy+A2Ob9v4m6sP4az471V/SuuN1qRmpoD+VsbX5kJMAghNfh9l1daFHLyN0zCyqcY8Zw+N0LqBOA
ClCS9Z84qMmiVwv/br6QV6z8W0YBddwKE48s1jzNCYGQleG6q+guVkEx3Fp/9qaNmgA6pYJbown/
J0l/0+24Y+aIxSaKM9ijhShd/n98dQ2mDFqBn9WrG6BcUH2xDk9uF3vh9jm8xjbGnKllY7+kVLCT
7yfasNUD9OChrZbo8NNzAo//p/DhpuLw403/Vw5ews3SVJ6kb/qUhmRghRqEG6rR+tIfKyW+cdA7
UfVduFcNxi/jK7xjAp5iqP9crxyJS2bIeNyYQ3dO9yKEdNdDEMcuLfTjNCQBZY1Q8+rjfPl0BNv1
YN5txoq7DHDVtOwMnHxh9Yw18828DEFeBomDPOBOrR7wU00pAicREaZ3GMsoRRp4CqJA4slTUD7+
ZNKU1me91Uj2BI0n1kSYTFD74rZQkz99Sg1B9Oglj876kbljoLmUatbYljr9/E8B0OJzzHY6R3XZ
dWRX5TxZ6578+VpiCVnJVp56pwUjoWDti9OGi2sYaG4XyKPK2GcKQSMfODiDU/y1+HHp6rz1P7K4
QAWcofUZPIX1GEXXDt9XfMFeEG7Q3pTL1sdzDDC65VTIMuCF9tPf8RJ7ZoPLIc7OhGQXPwyLV/eV
MoLNhoBkfL2HWac9437ge+DdBr2XiilAc7p8vBsd92Pb5k/Ya/2wBDyUD11cdjwp9czZp9acs1sh
mhexlxuFnWK8o9rUaXGRPfOp5VEUln6Ct2LbkFB8SnFOpE8xcRXxVGxHDL6DE/q+QN7uMk9RJGqL
E6ku5oyjlfa8t46y/rpjUOkgfat/40h/gmix0FUDvwx3Jq/taLKtoJZVh2ZckhSFYIQmCRFuU6yb
2ct+0V13FqBUy1wutgmrNULGV4eV79sF1yfLi23szJB7/fPgDW9jvBPJbIz6GX6eWJS6fImRmEV8
U6VhUADPmeI0V1+2S8pGRBSC2psYqc4F4m+V+6/RUYAAehchzwU2UOtG3M56sO/XSH7J7rZW+bvy
sFIXlCvRLHaS+ACrKLL8Ba93cxHDe5KBYz9X4KinhtOfe/rbgjvqHGND8qKVCnQ83bqCJ2oN+zKN
KSF/TFoIQkyxdjxceL5MWMsrbpEH4zK9orRqkL5HHc4Q/EEx09k2iYnLi+XxmB0yJ3sAKQag9paH
Us9BtwA72EWta5hwNAKKlHWbb21InGx+wsvw/AgS/DyJ/KszzQAnixOlFtxB6x1HIgFol+CnUE9T
8c03GWCknU7y5lmvHMDImXZ7pXXmh83cKmm9Fp1ObNpi1PGim1F5lxtwS0/rOjLvvL9aVr1Jka2u
q+ylnRA/HBTU6pCP5z8t6x8T05cWpv9/UIVCkfFgyL62iiRtxxtwTdRqQMO2MGNNfOvXADEXrBHm
KXq2ClZeeDq2e3cq3kQCfmKVK7+QOSBpWpdN3ZwG4m9v86JeV5jOWFYlYfcMc8FASm87WtZJHGlP
WkPKVMY01aPpp0PvwBve8WdNLG12AAeVpmgTcpB41MHs+HY6QXyivlMKl56AxGU0BX/4erQwq2Vo
X38feGokFpltz3tShZo/cgmX2TBuuzdL6MScvKnCm0l2IHgoT47tuDancgA01/hajftojk5l7geW
VeC/f9WGB6PX3FgIJ5olztamN9eex/f3TewqBXRgLJK+LX6iOJxVygH+fgCH91quoOIEEzK2xrEf
nhJLdi/4M7xR5qX86RxykPJ9XTdZu4N7fxMDAEyXursGV6leaf7ZW6J9NFHGc8hBLM6p+3H3/if+
PfmwCrXgDoPSvubxg8tpOXSlpSaCsyxyl6Ey3F8Q/umO79NZSKhKIMR8orgSmCms/Nu8TqKLqr6K
9+Z46P9GJgS1lbyo/9kcg1kvTDnc/YQAcsCjjO8XuLgJ8qYuebC6rr6maURVP9zckraJQIvlsryr
bIZHtHgdceiV+pYKTmAWTITsotX58gp7pWPrIvmCasdJXELPcw+kVfWkt3ttnAwoHXsDLqhRy9EE
V2rsgnsJsSXucHKCvlK4dfkwAO6cRus6vHuq0jWuwSQCK2kev26BE6G7T50BaI9hUKVokW5nNnK3
n4G2fSLSWdJYewGbC4V9l4faGGqAP3YXx0hJ0OK9opsikEFkt829LjEKVrHIBKpSNa9v6Ly0ZacJ
LGqAL/ujKvKZ3vvt7QZ/gKR2PJacaPpYWsXLjPvWFEQMHoz4pwGG2unn2nkBfLXkmUkBb8d3HUya
fcY1Rd7qUjTi46ZP+Z/4LnavZWDs6mk6fM/fLq9ESiKGiBbxd/B24Bx0G2qKjz82HZxgLjaTcEhy
FLPnJw9ua7Vs+SVref+fIw7xEQw0Om8IYf17Ry0CgFfcyU3jxg2n6A3iRBIJtULKk5GOtlEvYMNk
AsYUBqZexZU3wLgO+lX5iYik2ua6905HQfHk4+HqxwWLI+gA4eGW4MFIvpxUcppXAmWc+Q4H2+O8
bXkOAbfYlMPZKjb3yQ1WyvW+ROxDAjHI36il7rwswtotWKfCN9GxSx4vpHB2NpAJstMHW/Iodjtn
t6Bh1giiULGzobQkDEmGpOJFbyoEEpleCf1VObRzB63Z1lP8sMm2cs3HOgzXQyz+zzWX4qQL9DXy
aIeYwCu/XMKJ+0+b8q/S6FS+gfQtI5y9ZRhUW1EsH1hJ3HZaODCgGwzorRxRRS8w9iUg6klCNtYV
+TGd5sEGsB6aYlOPoB9agr9ExEcKPa0aDHAzlih2Tn6zfhHweqBn+IRSysvTmwUMJ1oKNUJ74vqI
bgjoZI2rvzgK+tjDLb/kkjAgLA0Tn1fK8H+ctO649T1zUQ52eN0V+CJ+0jE6XEsnyMFBiwlVJIKv
4FXG15GX+8FMlSkkch3ylXifSF3WKOH5MCu5IGn2x77BYiSyMKz80ZZF6dfrfIGtZPXlCpEbUq6f
psHw5ACqW27BGBPNtNWxEv93xfmoPuud8DdxM1qxBA5+f6e8ATyLMpLjkfyvCPi+ughsmjf8MrHc
gSv3NJUqf8rnwU4UxtwiMLqCtHS/UrsjGcxBDdxNNs47fQyS8A57wo8k2JcWSOazjw11DrevMGlN
KLdCn1yw0IcBL27LjMvDO0aJalIVxaP4CY0YWqmAUuBydSHiq4//Tl82017D2WojAoXxnjwxwtEw
IgfGpr72ICl7lPMg9l+j7el63E/yU/a3gN3UxZS/SUqZr/2KvZrjGLJPK2uZPiXar8FnYa72qTHR
QMmE/hm566CoDGWfTxfSOf4F29gwmj45XuQYuBlzsshZLO3tLX8zWIXyaylyvUtWSOUoHElOeKVH
k0XFTXNq0OKNZx+iX32qeTI9QlazgMMCRCP/S+B4PfExhEh48VeQwV+pNypASAZ+nProqRrfvsaY
yKIesp6fHKw4+PO5Rjj69HpsJ/GidDMdk3uY6t4RvsGMbCWEHB+TqOj1hLyPVsWI8zhAm5wr+Y6A
aferuYTt20gOZGIRqza8DI8qzWxGYUYUfiDD3dSqNlS62zJ97PF0bfrO5waHMAyHmGI5ydSDa7Fv
3jIlaFlPiLgfo/V4/YUJkSodEUN2xFHPvCzaFUWE9Un68U520uSpbHSsIHUFKAIeklqzxd+Syi8Z
E5FSxavod7RHOUxTLQLUJd69fAZirYdVZr8PNag5UfanFRn7KNraIeGIw2Xzsfm/JSv7utnR3Ul+
zumxYIiEkVHXTcig9SdCgymDVqj9z5UPO2J77uPRxj79VNrIcJCdmpuMWnqFbqRfp/ZTBuy8STTT
Sd1kNHJGNxYmVfi0lKQsXxvYtqgryzTDGpunHEj6o6QcVUheWP6iIaDMay0HKvYJKsJx7TwDUGrJ
Hveqzx00DeDpF/fgql8ltb+rpb4r+SzKjGHh64KmBKZs+pzZKjpnRuc5a3s09GjZGk5CZ6nbj2eC
bd9pl6LZ4K2uiNcUZ90rsVSfiSz6MGOt9iHy+u9RLfBF6+Ow08CXxcZpcv1r8BnpTrH3yYAFScuJ
Kdgg2HwWAUt8dtClDeBazvq7I03MIOol7zUQ4Vmx2Tajc6TfVPpJBcqrGFDzAN9nUgnHKXrthtr6
UFMVZrBOECz6eJWK/bS89QxuKnjieMbuA8cFNNW4URJ+PcV/UcKEV3Nmd4aMGAVXs49xEatTYNn4
HEZoNlFruoKncQ8MefXX0+2Tm/WpGLQZjh1wLnOkTz9V8605tOl0C/HvZtASBPKrI8j2PdMYa6tk
9WDyuc58Jd/o+JpUX8V381aHFW4ZfgRKwRMiQueGLO2wrOcE44yqTbUEjyAHFRjhVE0RdTZDE2eD
wHZS1NTj4P2MBs2CZJQwbQpu2tgC9Mk+LK1zo/hgD/a3lYXYusaF4GI8hw9P3pOEeHRDjDu4u8eV
JhqRqbJBmqgvYLEjHOvcsPfjZOuBdhsjQe54I0JV+JCdXDdI+hjrtuLIGmbWzecSt2D3+uQDJEpI
/xeQ9eZEL88xhwQAhBH5vb/FeM4KdAJuY6szZ7eVIbLV8s7fngo0CeyUti4RfPJVhgXg7Os9fzbZ
8YNRS3cIOMLi/gcNrqEgUynDtl+NhUlDfewIf6AW/MVAufYpjsNtWJ+PtKjaMnWx5sqvUIIBKWmN
qjwHAMTPNhZC8UK2NnS5kCJuO8lrKjnPEkL2wK5CA5J4QLRBGnZ00Gw72WVxq5vM5lZWDZ7/edRa
Chqz+S3yPJqbk8EzezHU1GFckiyKx7OVMMpqfpm8s5taxIeoi0svv7lILzzdmHGmWxllvv57vR/w
6lwxxeWrV1U4ipzIR07hKVJC0nqxHF5djmRf/iyuCpt5LMv93PPXBlrazb3MfxiU4nGBBqP3Dhhw
jo1gBJZ40AJtawug0am1w+0cRLKKNS8Up3bRckxLp1MRajNBh/gpfmI/tDBkJH5MS3WhwBdiIe0g
XqD5x/64vsYYsDDQGnFMxMiTAZlssqMIkdVlxCyJG7y5mi8yGPzfwr5ioXdl8ah829SW/mM0Mw4j
pILtbuMFgl5LEFNf39TmEiWU4AR/eDUQVY+LWPuiK+m/5JINlt9BeqMs+PZVnbss+AZCTkIiQiNb
9D/x265XExD0GSuZH+rlTCK1xiyWzD417LlWnXl3Yqr3Fe+ZFFpJhCm057ZT8k2KpXz7yZIVtLk6
R2+JQEaa2zHTRzc2po4pJ0c78LcDQ0MZRTJ4Jm83g/w99Q/LoqWrcnl7ag5JQqwvitareyFvEW0Y
r6xDYVlvaEz8eaB15HAm7EUuVQklpWes6BVsgYPIxkv0aHL/ps0WNOZgmrAIl+Iv4Yj9tTX9KNMf
akyi+lLK21dlWU2WgpvLdEZeeCWuwZXnCCsT4onB6T9z1W1z9wJPoBso/ELySlDqC9yve9UCIPRu
19Ggj44Qd9cuBQI5haa8uguPwqfbeYQSRdktCWWdkVbQxA/G/CsUxP3kT5G2DcTJrC2NaYT62wK+
yVSrB170AWo48NIrswyLRBHZEeJ9XQbCdvswVHcHrUpzmiUpVenGtGnfuHE7PKpN/s91p+6BHWjx
yq4C7RNBd1dRRJj1tARDYR/YIiB6DTOkpUXqWaHZZ9KVuPchNtJWuPqkE3mWIvy1wWZoDnbVfPkW
ZvYsgUNKb5PvFKFNGfBbXOAa9OrbsdGMMuyoX97T5T3MjKsocgv5ejQygo2rXTdCES2K4r/0dLEL
S6pUDkWgUzETevoUkCrupWTBsm1HGF9b7SKoldLPNNdcMVg5wAEtnC8vlBby3c978E0Sq8+iGexy
K0GjP1VVTgD7Aorq4iEQ9bhpulyhUFJMYa+vAfYynuGxM9alMR6p/ckVLd8p+5dpn/dF64G/wyz5
4g93nrrnDOcN1b4onmeYS10PTL5CYgQz7jMi7KgkIQNJbuPK/EY2tjKrJUmoSRGfPdTrJgZXEEQ3
tfY/R4aJSLG4XOUJTCJJ8GSXHfnMtRoOf7wSK/cFM5U0jmZ8+uKIkQrDHy4STiSxfsxmla2tJCNI
bX7Ia7j42ITTVq+a8B+Fz+3YwHJTkjBNrd02mlpmBjD2fKUqZI4AU0qzsE51FGxlbH29GoYCESKm
zpNyIa0IlW8xYUIiOTgCZUZnFw1zxnPFxN6/ZH2kmwjX4kheRUcJov1CF1Y1kN+P0ioJmt0BwhTE
04NSN0zqht/DUPqQCNB0u0/xE5UZhGQkcuOwjQ8H/9qNQl8jpSp9m8aspLUobd1ly/bCox6F/MWz
vfFB9KKdDwgjO9jMUH3rwNgSnwR6NBY9xMT8NO7/0r+RusBj7JqC2FZlSwQNm4ZYQWY87adlMLCS
dCkAbVYCS6m1EK20TSGAczXDbqijbR0/mu5Bj3h9JIQeYiR3ypUXDTf+hD3ScbJfNqqdKuqJItXL
hoIVOyklT0VxLMucAi+pgcIeXqdiqVrh0lu4ud21lolCU/XqgZf+0wEBBa+B5/kn56tB9xH14Ye6
fQ3yMoVcF+dD8p0V/J29qz+4SWkyHl01VbQWXrHKBztYQ4H8RPOQU8mpdapd5xLtcru4H/nR8BL+
+L3NRu2z2p05nrbGzSvlU0ogWrIetw/A0PopKDQBZV1AUf5RR2QLb57yIJFXiVO1GgUpDHlNFbPT
oF6hUg0wN3nuqYwNr5D5yF1KmdtLTQQ8/29Y9OP/W3DV5nK4oJle74XsCw8iLlahN8VwBFwtt6PS
GJ+CMbG5q8ZxbWrpCRSX+6p+HKpO5lDzDoL+zy5IJCQch0ZoO5zGRbcZvM8qyVvxERDNgVECMB8X
V6UxbxDrJtgt+cSax1MFT1nvaICUBjLBK+XCb3w8vOICHU+pccVdC4bTBvBa8897vxLI14Tf0cve
9eDAfbnyjRetBrFeRH+PWydlCqHpEJaneeGmtOps6sWTL3y6WkQHHH6CD3vmquVJG1U83yu1/InT
1v/HEtqPBP2Ybj4+BoN1JEsFIwu5qQKLpopMC6rDSCnL4eZOuMlG6YIvSsAaPITOYKPvaG9dG+og
7ue20+YsQLvSRhNt4bsFbFrJS7VP/iaId9zYT7kMXWTgIAEHncbQwU7+nS5mdfjOkDKDH8eDM7cD
4N64MTopbt9P3Y+5PqAyVicOE5lPsE3KBx7jXy9DwXmd1OzMGVVqABdU8yqCVT4HvBlNhb0ER3us
LThSUVwedK7aEa4xDhFHWeNWG4L6+BMEAbY6xU2IcC5YlDPS6lgBYvGfa6hsncK5VOT8RWaX+Rz8
2J+nhcmayZ6RFB5tPO+UlnObyPsX14fdNgnFCHrau0Ejo5UFP1j5pqgZiXsOdgK3aQBYTU8p1xj/
SEUqX/3q62SZqaLWOwD87hKo8+gptZ/toaofuCuz4GA70qL9eBNV/ZrN/DYafu2b1kBWBLrPF6S9
hleMW31/yQJkIaEwYmw3C7OfjT67ZN9lSnV4ZEumD+zfeHbmkub6TO40K/BFbCXia27pnMUh1kad
PzHUsCGJXvBNTm5dzKKaa4Hmh+dK35dZkIbujyhmYYl6y3ez+djkv73Uto99CUWjo9qKDhLVTd0u
J0p1T+eCx3fwrbaIM7Gp5tQkzRzcUfMdPger8VfHpZoflmmTYA32e9slB19z5DH8vFveF7pyLbJt
KaGPtfczdCpHIwMahJ2taR6WTORKrcb6VE9UA6s88AXyDm1fKXKOuq499DSWhHcnBadfwMc9dmzC
M0nu73/mtu3kxUT4iUJMP1ymolSEavWzCxvxU0s+8C+b4zbR7jT2w/4590OSa5HW5jfb+uXrMJQQ
tVv2774qRxGp2midQdMsSRvNFb35w4c/R6c6ZLkEWQZ2pJ3guqk5hbJkr4s8t6C+Ecbhy22WgPJr
pOc1IZgjRpQ9byD1jyKKzl3BMhf49yPyhCzSVNPZx2VncX5URb+hk8mWUANyeet7Z1JWBSnrRwZH
z+5/0LxZME7RN1CjQYhYwSvtj+HTNV3mT4XmLx3F9IeF3TwRDGb4D454PZVkoo/qMSe4xWBXQ3G5
NN6wgv5w3mubsXZtj7pJ+EfL40WlEm+ZCQb/aUBrKklnXgV+1s0xJ7D1L2c5fFkblaLZRGnviZCD
N6qUMVaFy8K7uEdExjgSjorY4b/BvAzMi/CD2/l5N8nKI2It3ihKPVtXVN0hkL8KwnXBP0kUPgT1
IlYZq7edczI3kAGruJm5pJ9EDd+lIPrZaAHOqilq0aYeSVmhvB5KJetqOkJvqaniCPXNLdLfQaGn
zlR00xjQ8CcZC8cNYKpIBWPShIXQBi/7ssWS8PkO1MdfAz9qKtHmqFXX+Qo0n74mdhnBQlruzmtT
6l5b/GEcmMZ1phfrg+jk3AI/r7740GEZ9YmmWY1/vlne6QW+eaD/850FKxHhymo4vIjNIZN70ErC
ZeKgS1i559cVnjAAq1WTXbgVihjQOAqGFSwW/YjSwNNU3gmeeanRM+d91Ek1GE3d8mqxOT7/MyqV
zq85SLZM8291rHM7i47UKNwfto7PcUGMFvDpXGvQ8sAIAbBQaToUQKmfrndb4bJ6xoHSBvjTO5yp
eRi4On4qeYWYdxY8XVS+VSSJMqgnzeEVtywhiwIFyMj84SPOKsPYHnHY6xAf3wZMOzbMEBHGC13k
TW8ARNL7tn0DUO1R/7OtjZAnhXOiwZ7kQIDECw3KkNY+/bGqyRyVsWerfpn4U/V+o3PlElaaP46q
Gp/xAcizDc9oHiJslvHAUFgymtFtMPkYMlGcm/6IB3t6px/MyXaZgknu+L4MKNkoqGkm3AQw/Inb
KgjKICf7gBsLjyvHWTO1jWa61yzfvU0IYWx4/BnH5EPdXww96Yh304X6U4vTc4/pNo8tDAlrelRJ
aRB7411RtJc0d7pZFsFvIS9ylSvGCELEfFxuRqgpvL1JH7BzOramv6GuAQVdJUZqN8T1/fPj8arh
8uEqNHWLBJNIPPib8+lexgBHW0KF82dWA+cq7xO8TNboLJOQMj4U8VGPmrRVC9NlamVLSOVHQ/Vn
8SgvIVDpi93XslvnXT0ojYYZaRGOo5Nke/BXfX6PXEcz+xan85KoNlk5iOmRmn7oVl5cO0XoD0Br
RWb8+WcrSdfqFFSZuwvG5ozCUAUtPgnfvMiEUwRwgILTDDMGcQmuoaYk4WGnaSm/xOTCceSuPnvM
fLdvFFc66HJ8D3IFionw8OJyZfROSi3vgNtXqPpYqRTEzgi6lmA1zTjnTxjEwtWie+KRFuiMB8c7
G2vmjFIEOFzBcJEg7JSn3sgDLd96z3jCOFgVdwrzRFSUrMYF35QqPKOEAIdX/Eh7b1HtaiwAUmP8
GA3PzNW9B5Zaw6WpoMkqrSpOA85k7gXSKna4/W7ABdyWf8m47X+xvADGWWnnN7/uyrKaorGAE0lN
bVh74eWS7rbOIo1n+f4iv/m2xus4/FzRYBMRim9TfY86HwEcreIo6WUPmcVjtT07p4zCUJsLmrS4
uXMncTcn6PbP+D3J9s4JU7SR6f58wp5ikBV33nwdHluN9OLjpl/TYmTuQgiBEZ18Zi31FjoUQYCL
dwRztgJPJgJlz83+genI9a0GZ3ceHnYQud/vHdxgot+wrZDgFrf7cRfuGfVzga3DRoVUGF0/LFun
FKguL1gCykrMvLlPoYqrRCz8JMJgDmQpB4yWuzxi22avd0qiLX5bw4il7exW1sAg2xUEX5/GVJjT
3hNg/FFec7dHa1GzEnh+1lu7apbiWPkivY1uXajC7GBbFMPWfJ22GTH9mUAnMI/Dgq0F3A106+HK
3hKffROr4wVR6zhNJZiJxLaDh3k6CcD+TpQRrDMgPJbTm/aUAiF6f75cK8Z+iMak67YP4FVznt0h
d9iPAO4GsnKYno0j+VP2mOqSAC7GnODmFRL9IT2Qggqw2yZuRgfCTQemFfZU3zxuI9QAbQDpFSNy
lwVIqfyG8hiq2+kanuzYpfAWcbDk/3DbLIjtGidd3MwRfprDcT+R+fwFG9UBzXuUYhWNmvbR8E4l
uB6EoNtBSKXB19RiYtNz+l7Tc5K9jJ9ObJOChwgctZQmhSMsZqBDVvFvFdzTbgq3a4+B+1BO7q35
6w1Q1ASbQCPNqVG7kO8Jd3P4uFBeHbMmdzP/eamxmfNyd1Za+y4jCtzLxRiB3bgIcv/ivCRPVl1R
4M42tBmzkjZu2MWhQOX3X/PEwlisJ0lT1bl5MRKrmuPgva0tCuEzECL0BStiHHmrLpWPSdIxaNBD
tLUfiVjGD6sFY/pfsTk/RqblANbtLrCk/V0UTC1nuWVkQh/DDFbI5jIKgvbTYV1h4pYQkrykz+Rz
pokTr9VXvFbVNhgEcXDEoRl3rFFEyOwXyswY2PEPP8NqJYmuQJBOwwS1Lrt2AFYlkSwOLj+1urh3
nKV1SdwiXyAirCpudSy5b6vzbojYPqWcDdiuH8Bq5+O/XVCrXpU3cjpvV95TeN5/yZHpM6RdLHFD
P8AN5Y9paCiRXjaIyw3zJLDaTCcTvVD1AhL70hEMGB+LCkPcpW05uWYVlOMuSKKyWJoFS4bI6S1l
NzY+fquohqbf4KDBDkDQueo85U3N8aAT0PZ8qfEV0IM8YU9BrFfFZm+oHiuQEYADO6GfxNYj3DJu
IHat6UPnvMDg3USbR2ZPU7N1d3vrK5EeUI2IlwBnCO/nuOBF6IJzaQ2x4aqVTN1tbWkB/lO27CUl
9gdQD68Ui/STYY7v4GXNptt5F05CDNqJQYfVT9Jt9vq3OzZ2llWF4f9d3XoSKc3UOHaEB/MpUNKU
73N8M7IMK+mz3pO3fX8uFQ7Yfdk6GUsom04wEKkLiOJUAt0Y3INbyzO2bX9xsSLruD5EROcfWVJm
bvyB0FEwc7aYT4i9RRdDms20YhQxZw7AAiBLZFGnBssapSbKddEkkGUYv+/9e8+A1e/zXGUgPYm0
oJeGkO3ogb+Gcb4sLXzseYtUmwMQ9AdpxG8FFXkKoxpFK0oOP+BECVxjPMZazqbU+CS03W584Puu
KJRtVlS1K3SOGzE2J/BWIa5RubQBhGOCXG01msd4YTRVw8PsPhozOkuuZpaCaGeX7+TvhK64r37/
NNTPasKOzndrU9dmP2UyIU4ijSCepNDaSE73eSXNi6pNgk2IrdBv2axVUwctRmbNqKSF+qkIBJgM
KtcHiAJdP5Zztqe2OGLxXZHiPCTJ/ow9lVeVwI0nz8JCzAkjj6cvfdRSDNXXwZ+UPusW2/H14K05
R4ahaxwIdwaR3MqHrICnNDIc/0Q/efdHfDaBMyvHt3lBZxfv33y/N23jJcybNIXGg01Qo19RMPMR
PBo4e+wVipg0GjA5Ov0ZcIMzNQGVQCz0jVvxUDcC6jNvDmRnW/XQ98xKI3jOTF8LeOwzgR8OxUwb
0ugB6x+XdncAaoxj2RwskdXjS75lcWm7vx11ZK5v1j7BK9wvo0MoBK2ZmhHrEl6v7gxcc/3g3jkB
L92WVobtjVPVVWIOtSEjKUXiasxxQMQL4UIQJfcB2st69SMedV7UULnewKq2Se4dyRcZm9McrI4e
DidDwDeNs02ZmpY4O7/OVauGnF2uRXQ3TcCrkP7B+tttYVh/RsCijkN37Fcw24mAkoL2/20Wi2gf
CJxQT94joH8Vbc/OxAYeRb7gHBUTbUyuZxw9TCt0e+VeKfytC1nn/gqi5iT2AWVO+1HhPj77BVh+
O7+veBP3oG2tOBlIMM2+zeYO2Md9RLaOyr7sED/P7YryeR/+lrOQM/7QKThYrBBnfHuFX5N75nZE
sehPH3hrc9JNl38JAB9L2iavsQGNwNcOvbR2ILiUtci2EX2/gV6GpZJY2CJLMQZJVj2GCHegycuf
BATbw+YSHR8BvpVllFqsav0OEI+cw9rv3LRmHgEIezk/cSn+qK+A9qXKXFpT1esWKKNzNNL9kNb0
92VsvIIw1nK1hENsJ07Jt4Anmm5OZGUgJbT2ulcnQlWLHYT2wPH1brAPSsxU6CJnEJK3T/iSgeHz
U89uD6q3INbx0LwysbXGU7j10NaGoGGPmBDCKg4RfzauNxOXSVqo7jbcuuqBRW4CcnDUYa8x0QrW
hiv24ESHVWElVT24+vatUSwyNRZj4OIWq8UJ4Y/ZWNQKz7hpoU3lG8inQSSUto4jKBCghuZTmJAG
WcZS0iokmKEsDioQS2rS3snCzbliF8ZHq07VxyqDJWIKuwZHFEQafp8VtluERyAbid/W+MW8MB7n
vM2fLUZN+fwGZdpdJwfIre3biflfXl+iJx04SQ2EEimKDtzlCImz7KzW5iQRu8BhN8WImxydkNU3
gTCUtMh0wM3HyisNKLITb7rI/yDq7Y/gqNeniptf6bwQEfTr3OejCViU1n3tSp9Sl+qi41owaKJG
Ge/R4g0VMoX15G8137EowuosGN0+Y7BUD8rlpkykug8bPh05nbcg76DcC8lsPha3ewRbooQmYERd
RQiSRx/zvwo9TGuyO13As2STTo2gsExth1mjSEQnLbmY4uhDFHt3laxE9R/yso1Axfzmjn5KYsH2
jLatxvbIVx8CMdRFXHKlM+P7v6+b+iii/IueWi0Prmsd9uK3wHdJUycRhqHBgY6APFKYioc2R0CP
V9TRWiS+oUPbMFUwEXphdA6qopyMUnh8bFCEmLNB3mXv+JcfsVGK1Trg54pcCHWtkHQ/iey7Bog1
6xSlfPI3CEZCWi4Nd5mS4Rd9FfGu2NKZ8/GvyVM0+AtYkkvdTlX7h8xp8YWXSD6zmMDMMLW3cSQ9
V1kNpt3AhiQ+HGFB4Ihkqq4E4uxQymT4sRNy7We/joU9Ek39ehq/mVE/oWpTR1Randu0N7rtqN39
TS2gHSgbpaE8vrPt6M+Q+56praY5O/gb13YSeBZo3D9XDZcTLXmtdJ+c+Dspv0YB9sUFdZha/FwR
xXHl5KeUffyZivZOwJ/ompnMiX5Krcq0O/+gcn62ZjzgmrH4x3wbG+xQvBvWkG7zyeTZGL+2yY8s
C3tNvuL0uXStqYOQvz1r+P+WklB4K9jvqj/4vP9xNcPpxwEOEkE7lRduFfcsYC1B2lJOS1Mer699
U0Zlc3zfkSau3AyqmsruLDL5ecXZsTuMXi9uzF8SUSOLkB2su1O8r0QuKxOFuAiFDHRs5rCkXVvW
L5eTy/+wAOrC51nGoj2ArCpAi6dYqkPfVEJ8WjfpIcnoQ08cxiFkleGuEge8EdkKjzqvgKYNZghq
4HNl2fAla2GS7RN7AEfNCr6PGBh2g0DkpcW3rQRGzFj7J+M+R5WXjM0tIEEMWJ29rC9J/Pqc8WFu
Z32vqxz7GFJ+ejCEr3p1AAOrBTrwqTgnZN3FuyZcDD92Ibo+iTIhG9/WmeAnXyl4lzQ9geGANAPT
/QKhAbKhbWqZBeS6y5rz8FPk4KePhXIW7n2ZxiKA7r0Yp+gXrb5gYVkFj66VsimJW2ur1CPZNokI
OUYDqUwDwg2w9nFmLbMYNr6dfQcvvnJo9n8r4p/cNy5zYFAS7cvacn7TTwlgFxB9n40ljx4TuCxt
FdkOu2872JxCMwjhveAvH/M+SUb9gdo1SZ2uqIj8UwfpnT+M7Smwuh0NE4n6hAInkHgJjtZSNgEV
MYj18W+SvDuMp8XfsSXgQACnlXm+2SnIoPrJxFJK50Lzx+Xku4lxk7UF8MMbWCCas/xkPYb0fC4c
JwiHrqS5vYNJp8AqolhY/3avunRU4AmOAT3uhBnWtHDSVl6QIkHGUSqByvqa8vQPBAgWNnav0IOv
5cs4kY6Jqwc5u25Y9d6GvTDQyBcfSYUlxbOKlQenzrzxnQJ5Iw/zbTrlcL5BikUjc5JM5sz79CXI
tiACIY4kLJvIYAkutP1h+G6tOhTG3StfwfKZvOrQYoipdtIZ7iL9Pw6mxkT/Q3+JeM/cYEaqzNkt
pKL+3jwQIjOkdAJPm8jrp9NcdffJEikRQcyTMIZP0eYRdzR0bugStTgwlvwHo/0zYVdafYZJE5yG
f5W4t/XflGXrP8O6acZkiv7jQku+rtUkpXFDzTsLkHFKLLdNDm38q5qM5VeH+Mm6d9IzgV6F7wFe
gkRHqdWSKVrv5ED/G0qp4HvLvlGAKQvN//E6pNPu2lgjfqTztMPfgW8qnpsQGZ0iO+T7Ue5lP02o
gbMxxWXBuh/7WRUiL4EiIefON8obB9lI6tuBbu2GAGUaKsBJZR2WDqDJfqO44te9oXEejyk9r6Qa
kfZCt2CtYiYzQ21YXDODA3ODEqqaXKFVcOHLkdtuegNEmaBc/iOldjbkiMC7DAe3b3nLyO1FfGll
LeO9rgy71kGU1mtxp+yIP9VERiLL15rJdJDTL7s/93hWHdPgCdTglZCoHj8PnFpWTLQlkEMaGxAS
P7jx8IA7UtPAEbXsyZknuPN374HqZ4l8nUgycMT8syHI8EU/dYlPjepd+WGG8REYgmVGdXu74Coo
XBshgdK7wd9wzWbmsLu/PK7miKd5BfDN6cVEZOzEDe+1qBLEl8PQ0eKlb92CT9U4zN+S4AMlWEdT
obh2wONZOtzlVdfCV3gqPJQZA+bDdyKRZSD02skfON/ScsgpHtqq+4Pk8haUJq0eJEoOO/Sv5Sqz
l4urmFAxxob0eTKQL4ARtJzxV/tUJT/JMFIu0W4kgDMuDhMrj4a1r4ezTQ3tnRARl6c8Y4777kdS
uvMed7Fo7+tn0Rd4ErELAc0PDYq2Pi0vFAtmp3Ko/QxaColbWA1WG5aq6Bz8M1XfHQfJrKvWke9B
m/1DGORcBPc9C4HpzxPEPemPoeYrLUIPd/P8+/tHy4kF3ESJPz/0KojlbUZ03pjqMyV4R2GbF2Mi
JFME6nrx0bZN3+4PIeWeYk+2JtDCKjRVmRRHLz+MJOaft6clu6oB+bXW6TqWeyMe+0a/Fc/HQqD0
Pbc4SFn6+QVvXw1oIPZz0bKLt1o7PlniBiG8beg9gMF80VUXlAdBSKsbIMD0aFJn2HnECQsf2eMx
Atrux+V/61PD9KNmF/9GvLOYGAIZFWNEqr5bKi356pj9Ksp0aV+QlrPqVJyZn6SMXGkx2qzPQqlW
Sz/nABK9VgN49dbUl4AnjEFPSq1phDVgJ/PwXLhcaS3X1N3aG0hCxEQMa5RhmzZGJnkhXvPm5ORP
Vg8y6LYSqrSgyTSple3fmu1Asoxbi9aklAyCcMSEDcawP4PqPtllrg/jRdOC2dLctxaMtxrU/AAV
S0K99/mfvJxfi2Wdp7Y+OPblQsi2HGxbDolJarBT3Rizv6kvsucZ5m1jQPrqCSyfru2trnO9tdgE
Tx4jMYh9jn7aDyCN5QozzSNPHQNvLp3UiNCCALhSgTCbhUCU1Bs28FxkmdtC31adgQHEeRZTrAFC
xG9oPWcpgmBwL8KdgeD8Dn68EzwaHpA7RIMXZybw8lp7Kwx7AQSA5yvNIUyRJ18CwlMYWqQTYnM2
7erbRKWys2m9qj0hMgNBDriEvmOWPJJc2Lq9ToXXJ52sJUlITxaPGOmRKEtVK6W2PziR6wredFGh
z9ejG3f4EGHTXGGoDxoSZEZY3yMjsvDksEr8ILxMA4RDwMR8Al+oyWgogaYSvmShaEQmVKTshJKg
gqGwHIWwQu9Yj7DnrfXTz0+MoIPYyvwfu6/FWbsLAn4pNTu4DVv4n0Q46I0iXRhs80Z4l/A55NmD
g2XzS4spkPp/+PsHX5dqKZ+NuaaR2j35fqxqXJjTSCFx3vDcQ47+x73nVoD4d5aRMxQwwny4cmat
U4ndz1vKmXArjxbXacUv0vExVEykAS3jIo+de9hy/5lJie2/6+IUHrAna3xeDMNfaA7JJkbZ9Jon
TJH8fBNzgNfxgJfEx02INlCU/S8rw3lnDzha66es4POlC2o1PRgQDtb7qvRbeoIagFaBPwWL3qB+
epmy3bA4Qcu/vWRIgAErU19HzPwnwU9hNhQ1ltPT9mfoMim4xb1mkz02jDAQSz8RD5uBWtc3SYtS
JSK7FWTdolQyMvVt2TJTHVL+sapgrrkADj357xTj0AvTYJ8UR2w7uN08Xqsv5BHhZ39PrTyb7G8g
pm0INM/+U5XPDhvPdg4Za9E36BBv2DMm3nkT/OZTJsF7ROZcOngcTqE4rZ5OjUrRo9E2Lap0ZfP5
e+1U5jhj2wnVHxpccLrZHtykcN0OQi9CLMs6JeGPLvoDtV7BPqBy8WfGYFCUe+X8bPaEIbylWa0J
MtX3vusIXM48HBlBZ+Ayo4SNbmUprQ7BTWbbLLv7cGkgIqrBleySDaxEd9cZ9a6ecFVFyASglH1v
G6KznH1QPs6pKWslQdqPNmk55orMgQUJ2X/aXIP6wpJ1gSbsx/vpJ9Do6pJGj+TIsyZBxRfAsVX4
KNqZkQXOZMGUEDYVt7cWHlL7eTszyXr8Mbi8pAqrm+CvL0DLwaKLEHLWXEJ5pWnb1xYJ6NzQbj6q
qUS33p85zNflZYsHIy6XTNYnpuJzgubyqm39Iq1+sIHtMqa5M2M0eVZwBosg9aSGR2M040O2JfBV
PEdirktvF4WoPyq99hTKfn+qtveCMZLV72xXDBUb7e96A1hcoI/dCFSopzBp29DFQRu250RBKLWe
ADUpmR4KoEs9YvyWx/TdpqJLWrTSMzywMML4ELpD3BbrzVKAhAD0mQHrclG9iVQ5YnHUEnAt7mxR
zb3CFq0w6LZruI1sJXUdEXnTtRLjuZVb1nUOZt4YHljJSRHPZgeiofcWhK8iq0YQVcqOGxCicNbi
NiI4SbLt8rJOspd+xZWB8xIfcGE07Fq7TVVnFPasR1QHhCW1zKn3kcrUiya+Imff/EWFwaiQJhLC
MuBV7Qwsp54bNyAvgTYcbWm0fUYx+0ZFOtzd3NZrRF+0lJCjJ5GFfFcdaeecECk5EJK+98AtnJjB
VeNCoZySJz5zHnu4YcTkTKPInP5YdY3DZUdRS8s208PK3OZ9f7UJbqGn42FwyDNJD2PkwTAXYY0D
xVRAfFygsW7ZPsGv6ETsb63IVf6jiHaBQZAaqVryVnOsljClAGLrQBMIPZLNdONSXR/VZql9y0hi
NtO5SLSrwgKzB8FovDqI7lkDOKrGwkXRmSQ2wBQ3So9MYQij+L62J3q+VVeg2UvEqBR5u5gCDgob
a+1rV+m+3YYg3yCkkG2KNHfXi4pcuG7N8Bie1Ey767hN7CqIlngOSD9pgxP+QHmgVkE2xOwsUCG0
9hemDRecua7cpLuYEv+RPWATgtzPsLwNJ1JCFWiDOd6jWffThqy8mbMj0vH0ytX/WY7FdfjEJyT2
MfVgCFPYdWyrirIJ/DjN2GuAy5L4jki1PtIpYgKG3JuDxwM9PWY7pyo5S7e9Wx1Od/DIJoClZCAW
Srd28TeALVqm8oK8TlmdrIWAiwVtCEeJvcxlXQWfICcvBXAEm1OLb9VBnmFVY4RTkVqqSXKfyISM
3MW6qtyxcFXzI2gz5hf2nHQ3r2vQhNkSAYbIdHhBgqlMPlxrcff+KjF5kHKG4hvNptEff7MF8kVb
K74xhHg9a2FEexs/kUnOOnTm2tgWsYXpFveUvJoAZ8AVCSuAq9eNPxvVn/pKZSfHT6dA8vDRNfVS
DfKABgKBKsQ93SdRF9YKDnXIbhg/9U/ydSjzGXLLADFH9Q+E0+4t5QhJBaMSjvP0xBOpBNxQDnHl
xNojwOhw4uQHbEswIlrM+NWGUNSCK2eTeo5T1Lm1a7cbJLg8ukw4KMieGWBMfc2YEMXTtT3IvTMF
ZSo6IjhJApLKGmKXseuMBCqJSjOSgnJ63yBDASq4RVrdYJR+NdSWm4s+kVKSICQDl3US0gGwFuUX
UWRz3Q2PawFtz/kAsHBBoXTeSa5yO+scV+VIbKh50gh6ptKPlXdsTNV0PQDq9zMVyN0kPsaJN3Fj
OErLBCsnnXmT3mlRjFT0kLKa7QM0lyH/Vt1gAhIT8EpLSgj9qFJthXZigZXjYDqYVck2X0ZlHjsb
HrBN0eWNP5HHgVm9m9e8aCG8lT1AiFn9+B6sPdHQxIp7QRC/z3iT6ueEr1a8xNGAwISrsfvpO8kD
GaKgP41DIvJ1gv1aZrHVJUjV2CENU9KawHexAfYAQ0NyYPBVLfAD9Lv9fpaFXp62FLTKckxFyGSb
iD5ldLQYth1MvFLkkSYekQZxK9PNYU3i/oxY4Np4Nd683Fi2PYTsZaPEOWH/QQ1flFCYtm+YsA+u
dSAJY1JjbEuNWup0F6cZOO3yPb+yn2OLey+oi1Tr30GCOLPccHtEHa3SNK7MUQFYlYeLGgZb51Sx
tZfl2qBji8A9KtLJeXwZVZzK7D6YkSWbE/OWDAkMHf7CJaCFsRxKge+x6au77fiITmTxGozzAvDz
XZLgW2faNhwYnXZDwuAond4MRnJMqen8YUIqJ/8wiwL70Gra5RR5ByD6v/5FBhbittm/vVSSp0zC
7uldeXRUP8L5J1FEXjyzyVUO8m5vM6UrtgaXBs/HNyc/q2BAjY/1ocq9Qc/YpEWFP6kxN7j5cYCU
x5bC4sjew73X8fScM5kofl/GZMbpiZeS7xRp69BzZNKs8AzCuS4ZkMKK/uyPbgmCALdzhB7tLhwx
w9bzGl/mitic7A/droBBNIptDW7W/vKyANj5EcXkqrtzZ+8hXx2LtfZnHY/pQBUhzyMsQIf/NIIM
rVMtL/SXs7idr/5I2sX18muRgLIzcodaRkZ2u/ZeCu4QE7/o+dkGlftEmcvn9RpHs+N0b3eQMCvB
1DJ9HDFAV04/Bufk6sc4u8TR05DIaGahbZMZuC5EcLnorSfRbonsZhCfRU50cJo3hPHyPjD1HMd6
DLzT9EzGWMHqgSKFFgUn/uF3UVCIG9y4RU1hAN0mqlUh6JndTFfwLjEhnwekErCceuZCpIdDBbv0
ouMwTzHzfotpu73wcEa5CAGJnjBW7z9lV4De7p0hdN1hh968GwgKLEXsQq0NAcw+Kc118alsWTMK
idbRj3oXtizhErhvKtGCOf8sle092OlgAOSkOI5uw7kwBlp43a9/G0un+NwRzSRrCQjbUSE66Utf
v4yiG0kBu5aKzpBsQ8tsuzwFK+dPHkqA+kwu3QtU8dWpxUrYB6lzCeMuky/kcUzjOvnlnS1xq4MJ
Q9rYHPGH5uuMtVD33fmY2bo//FzgArBopGAd3CdSvcAj1VAHpfmUGrEGF3HuwjzxtuEibxt5g0S3
7c0cpwoC0UIThXOnrCbSQbEBTNjgD/vc0RWoT7YiqLFbwTiAm/qOdNvi32SL9KysR0hkTRJa7JhT
Lph97smOWdT7XTzAVQFK5mggzzSycMguxvFfqgNPsN7oTeEDhhbbLFQGoU8PeLgjdRMZGfdUjJA8
exOQIyrLyDalHp2mNDKtBDg8MAEl4awjJTUGtnCfLAXU1jlTgvPDy6tV2mQPaDxai1zB3Aj1QFrz
KnRkd6kmaLbyUT7nz4Tz9wdgGDBNo5YelGqiE9e7XBUVHDkIxmYsUe6ugqCs6/tSFwW+bdtdacLG
8TY6aH+kyDsTQ1kASkhKAdNgABMCAOmeM47KFXQbJ0AZLMTtwc+pN5i/8MxdkMY1xy/WRJh6rAB7
Gx32p19PYldHw3y8n5+kGbwJTCDMrsfvTY3i8zQVwHgi1OTRGo+pJogodoiZbV1Ep5FaCls4pkv7
GnRHi5eKHB4RKJrZieQaOw9tbJ1cnGq2+91jkvdUWLVELGC3DgL9mceAJJIGU+OUXhIZZsgGODcK
LV42UVm8ZM3PEtcl1wmqbrnN8A59FirMICQdEddSoEioGS2kU1BTeoJbjpMJZncAhum2DwjOdcnN
QjnBaf1dkf9sGjgLEZGEG4Z3+KWrOGSvx9x1OSyMWrlwdGNsI9xiIp1bG7JwT3jZ/d40Gk3MfFbC
sYPd3fecQ+fBmR0/wvnNOAWZIHOwcg/lxZz8tL0+bL77vQxauZKesxjkO4EkxxZG1l+RT453ABhO
wQeU+xAZRrGSJGnppESKT52INj58mKYRPUwSdq8b5zU4K0JI4v1w1+U9vx6s5Yf/JLs2BJAfXXEd
q2tIi4y4i5Tk9Acaty7Il5iFMsqw4J9ZFfQzjdyLm5vbAG+bjDktKVLSmhTRF0nTMPcMbB6/Ip+q
G7QQYHgSfw2aoMjgcpX1oT4xax6UpDzQPxsh7nh+JxRKFb60TgoJBEK/31bH8hpCQboDVTMrLdkc
gJy7AIljNnIwO1ZVGk2SSmVaa6zcMC7/0UqzInkexriS4jhDP77WyAWJjN2gy1VzLYEqsjZnvcis
DM/DhKzjMDeV+4Wco4VCPUsioysQ/VuDrFVwVLgGwbc09B5RfhmeNwtoA3nSy76yIWnzunIkLpyz
g9ayDFiZle9w9TM2EbuOLjmlUgF6+kMtKfzqld4tQJ4mY0yNFQsSWaSIKKDwvCrszjffkXtBD4P/
uhFZcfu8zt1251FBZF/rAJKoN5Wgt35USPQpcHnyj9OJeTVKRElmfKmqwCNQ6ykuDEh3I1/KNe+J
mVcq8dIuwWfN5kCFsqpSQwt9N/gAjknhdbelY/bWgp/4H5OjKmrKCk1HQaxT8j/YaHX4jRZvjbPt
SRgqVm7rnJhLqZIujt6uK8B7WV/CN/8E+8kGiZCMsHaNN5ISCuvSytfJ4nB+R25b3qqAlH5a2crs
mgZTdBp+dk36wjLDIsW/PiRaoiiYV907P0oYCigj9z4K+0IDvLjOEmLnz90nSlKY6njuaFXgo2IE
QYol6HjAoTGwwY92dN86DcWQ1QG389qxdCcaDG4rmdte9Am9CXHAib0RgiYqIKiFdZMNb9F6yVeg
+fYcusRqMJ8WyVemDIUkFwcWfd1wxdw/RbNKKiaQNLV1AVqH1OuZdf4mCULBpqw/83tNHzvXZuvu
7Pfi4BegZhEubVD1iFwHveZ2YKvlsQeHZfXbP+ghkX013ljfes1lG3ynddpp4c0GMrhQvC2ix+sg
F/FBiHIAcTp49wfm6nwEuGfm5aM+TdCDqo751PuDV71NLjsZMeX9jjOprGINnpHCSXv2WfPffZTa
KLBW2YOLDa3TLUln8YL2HmulSZte5kHcEfybrrNcTAucR5mIZHXdMYdmvcPfsPcgpCCKWJDBRHWb
sFrBV6GM9l+kC1o2CNWAewtPAiQVGaRAxL1B+ngjcbXXWF5j43wClhRI0XchnmAP9ImyzkNbMDOZ
DwAW6RNdiWtOSh3eju8XRvx88ShfgjHJ81p6UgKNhdqAaZVtZ2a407ll8dSd5VmKPGX5ZKIKg5ts
370CXvczrXWdTotRZDrv1NocN9FvYhVuoq4/oQBMayBEBufJiBvPMPrViabkzXbXgoJ/DmhcAbdq
jKCXvNbARaVPCyAWUMqT2xGRgphEEoxk4AUlaI18utfu5om32qq0B3PaaEVedzvWVGpZUDqgazln
4YE53OxtPW7RMoFbB2M2W2YJliWgSTNYnTUc2OMgjd/OH+aMiKKF6BLu1OzzryvIw413cNH6dlVG
UKuVupx5Ho0wTorzg6KdloemxX1cwMZXRC/BRceHzvNalEhRr1UBoVTxhrfFujTQIcrLrkLBLH7M
pn8LCtgeoUrsSCXpixtd3r32HhtDXDFTWwgVgDQyKClJLL7A2RgoL6DxgqCqJsSDwks1EeB1+CSa
0uMInCJ15MTI7rR9HQLnowYKCALWejrhsLsV1mON+DBF6GfT86kBEdhx44Q8yL8Q+SG00BzWHt0x
gqXTos7HlfF35h+D95M6A19IaZVjAUP+63ynNMA0qb9aEMCXMssYupF6cXft4/CnAOvhXbTgEMvM
lSEnPSpcZQsI73PnLcFco+WfE4zL1MWsrpPgX3EzpZMcStCnZ44PlooSq24MWbwb6Y6VGtw2iqc+
A6ym4wClXhwnICjTVeitwZFclk9cRcUXujF0VFSkm/7YVfAqI9bC+xwkFe2XOIHM792B+goR2KvO
afFaM/zsgohVCh7Aq/QAtZ6ajFCeUdd4F/Tv738y61TdoUANK46wqB5ujkg1i0y80rmUdfZp+Mg5
uvBhprmbGlbrvPMwRBv9GZa60EHjS6z/c6pNx2lKRwo3AkuA7ZvOJmXwLPWMfFHrLJJsDDobiArY
EICCEnQr/OwvfVdofEEgfkLVcNtu4/FZCzmohAN+szRUHuJi6wNi7C4jwIwMGYbUB8ZZp28zVSR+
mOOy8Ht3/tx3zORPGxvVkj3tFoUfhyBP7Wtc0MztWLV8xQ8CfIWbfFoemtSFSUyUhuUwUio1DeNi
FS1S+/blSfw/iNffpQsCKnA0ud5ZnFIvIgwCToeA0ZVgErkakutpNto4o7jk7KwGGfvrcVfJPZIB
XPoKibK9Z5gy/5vobPSYzOiBNjQk9SR09sPqt15IDuttc5eOjid/aFWBeYwSx2e/XmL25Fnu04Wk
pzvfjls48Ig/OBtacEordYeV0DRHRRvczQVH1hIfZ1EqQNeGgJKoLfdaejEkrJtgj+FZgtNftujF
VuTSZvgQad8+kCpDUPjhIWZ4iHfRYQDEJpfIt7qYe2gsRaDlhIr5NFQWHwLdUV8P8YVRid1r0IQD
2rP1cbN2HJlOO6Nwlk42Y/vqnpdcaSQs1QceAVRStSSARxJrlHY8O8WoKrC7Ib8nT3NwUDYDUD/y
lKMMeOrCuStGVPh/OFAgpWhv4E9QqEe2eBQ0veV1t78FklXYs0nS8b1+43HKaDVVkgpGe5IlZCTB
APwhOkRRqaBizSq5qV/Oq2fxPbbFcx/Sj1Pr+TFo+bhu5Cj1w03l6EWL3NisCUoMxtQ1hGuulRc1
IkQ9DFAazb6INjyMKFU1R2qhZymRsLuMcYQTq1LuNjQrXiuEL3KM2raz95seHWigzKhKfrw+MLkl
2W7gXWMVls8Rl5XCFy7KuI1VRjJ6CoHHKI8xA5OVDmFkUYcm/JVgmnHb8CYqEKtCVr9UZnaYPnPH
OPtH4Lx/NFe++IvB2bBqa9RsobN04PINIjURojwd4dePiPZEialEGZ+oC4J67q/iasLrcXZz7FFK
D8uascPqyGFbwEk53jMQKjgjSvHPlgV6RTPSe73zgG9CYk3enpKNxYm6mxtJhXf02RWNlplNAtOV
uSiY6lxLBZUWaKiAUWCXJHJmUM0nr9JUxI81JaRQHQLgXAbZQVm+FOF5ipfpB/z9iSwV9+ubYP2H
wwShwdm+z2ffOzhcHvednITeB43rMQ78k3p1p69630epwYqf8tD1el95HTct/+9w+SRu5qpDfLTA
pkFTEJpP0ssVgBqDmKShRDI64w05d5EIbmdJhED1TdhvtNp9G5ydtMZQ/vbPUcpMP8surGCHj3qJ
1gVfRWD7+8c7cQRbJ4eD7zLg37QZGynHhC1QyH9Za+MVc5wnYOa+qPYlID5NhsR7UGAPcvC6KzmE
CAXF5nI4bEtszFtyH8DMsd+DiB1lKYj1btBVb6Mu6P9UUZkcYNv7u/2nFg8gyWwa0we//3GbTEp7
meRxu8slKREKJRIjqvwdJj+tUciUxBQCahngfBovozDfxUYtgu4lvFYWtJG+urDl+FiY0OqMskqL
/4xPve17CdAqIxD90AAYKIFh65Py/6kbyhYA45CwVGfy+YKnVlnxt93KtqmRw+tyUrf7fuS8zCGq
D9hlxZuDDb2wJY0v7Og2cm2wWMj8s/KiC4T2/poD/esOaOEbu45cYvoccbyOBDiR6zu+Yxeiejfo
+wD2nxevck9Dy8rZNE/Eag9BfEh2wD0r48jAr+Au2o/+zrNcbPOsZGflO3bwbWeBtwwyA+uYlwcF
XEN04/tqzygLPhpi/Tjs1a6hLDOeZ9OkPPhJk+eOzLzqBXOprIeob2bui/PFbOY7RarJQCohixSM
eAwLzKiWFXefI5+wkNBEpG9uJkD6WUB7EH5n/NAJsiGDbXaSOsN9vM5QdSa9VLmXIZuT+TMCgBcv
jJRjvFPC0mQ+W/46d2lhA3hxE5KOnNIOk/qTM5uE4lwyFxOjDmsnDOg5/O+ALOSGazOE/3881DWf
iSgZRe2u07GS+qMn0sVDNOq5QlSGIWZu160UNHjc0sBI/2YjOi0j0ZwVDMpBP9sOdU9MzkEYcinK
mfp/cpVJGcVJQQz5rgJwHpcM8gXBsA8J12lwI+Kqtv2qri4aNIJ4wGgU3GEPJifbsALyP7fQuwf9
iZF6PBKDONUrviXl6z7BY4/OS8aZr/8n5pEgqQPYCH1dmuJmrqgBr3jPIUwwBhlH7Fjnshw3UIjv
MaZuVomQ6OlBPlXtxlXDhTAJV+27ycVPWHeKzrngkJACKSooTV+s2U/JDP0fXXJ5u7NiB5mDgJqK
ffW7HTtMRNJlOfndMfBbW/4qlZeyiz2owKcxiMTlA+fGD4B8W2rmYbKfjqgKpxkJJvyNMyXjW2lH
WMEdd8PtIv9H6N4cckEUxSUZ9pbyCpNFsYC/xX2wk0iyzauwr3tY/pI5YFSArO8ygVvqjZ0WMssI
EImHvb91V2Hg8bonJSGplwvBGiEHvV1za33F3GjastZWYa1wbiPe3cbBGp0sgCJj2lM8X4Ka+dV+
ww2hrnSwuBpq/iRid4RYxSUheUY2E/3cKVCz4jv2WGSbxLEULUCBrgFKdYJ1lkE3FpDDIOsaBu7a
vEyiMjt/wgQvBMBSZCZ5clCcppEH72dAMafcf8GNgF4PKQOyMaTwxDtLU+NOBxtZY3TlD875SYKE
/YKd1ArhceeGyEgRWrDLYMfPDQJN/cPbfC+D9SxR+NFVqX7997qBXaxqV+ZjitiEYUwdEwUrBj51
OwTgWHji3sCjGOUmsg+7TtDQzKGw0JeCvx+DBajvakh3g1ib078m9RE9guXtJ3tMj4VgZGAbi8ip
P1PY/BrLDsL4x2qj6IsfqVT/UVyv21GkKJjQ0qQrzV3Z9dLkBkcx+3vHus5bOl4j1zpG6eL+EsoP
N95quhtOTCIYI2wxJdMnTdktH/IWHfSgfmjJM0bjLQxestvUTrJfb6zDQw6EuVd68DfmUUyfyvyw
/xggliiBl0u7fyoRXEuXVonLYU2+zxUfhxXNFmeNdYLbXo2zWcuQBgDnL5I9XFHMwA1HffxZTuqd
fChekIqP6iaCqiJa7U5pffP1mzzTKGtjItefUMHLtDVR9/rnjDLNWNuvLc3Llcrh0yEFyF6DMi/L
yOzjXdVqKtgykIHwsDIF99OlMbXWwWG2ahA33mF5htmpFYJ2NaJK2ZU7zmTA/7/dBGscuiJVRDlV
BoP6b0G6pRoXuAVN5fGlpkGWhNKpeh7HrBIJ8WpcymaeylqNLswvfujd0wN4mvtzLd9+1SVwt69n
Go9jHDy92NB2qmcXeGS0xFyyrVz2TTVrtuCSoWT4E8WVP2jT8177IpKV1vMY3ONPtPsYGa8Gr1rw
Y25rxjxBADHRO3a/FDIkePLOStrNrpBZjHZPE9aNLVKL+lHT91yDAT5kgqxdKsT0z558dnLrRsAG
TZ4iUhTt6B+olCeYvq3SbU8bmdUu4Arg/26EhaGNL1dOXTV+BkwktprxLT072gH22R4OLj7AoaFi
dA+DSt0PubQVQ78KNZ1GFsK2rAZcGPgCbss/w5xiwzdtnDrbUrjFYZdVtCPGUYLaHAnYOnobg/QD
RaW1eBVLz1vPZD1yFWuH8tiOY8osk0GW4tlZi2Pm25/EXhDtSEprcVGblCxo77agtFNU7K3gzEBQ
IPAxytbFLD8jlPv9l7dxgluTe+7LPbaxY1qudPKFPbS9NexQyfFr0xK+N4s2q0pPkiS1E+UG2EKa
Tlv81/fwthzCifQ7tjZ0o3V/cef7wBcHr+L2XqfFf7m0IziarXkGn7O+MYxXECZjAJfn75xub+9w
kajUg66ntVz2mc/9UVi81sdnwFbpkCNAe7pg4oRYNi3iW5dLH/FarODl5bEFHbtSqa0S/sSX+uk9
HoubI79YYjbXQ9sJzwLSymqbFOYdqQXZh0/K/1ivJVvw0jwWuXy+ptxRLF0B0cIVui0mhVifsiuT
OxpCSdqxn42zqUyuUCqgMOv49FuiQvdGxfotDdFRV1tIsoMMl9p6EfzHPPvI65SQB09yhynVDS4o
Ty/yVO0QLjmybl9x9jfh+mxPgpP+Ph0yOfroKLaEsQsglJgXI0ETZLGOpAW3hBl7kdEGQcPOFzdL
jxskYsj/qlMZork+u69GU2sTiz9k1LLux9mlpCoRJTEYpWg6Wq8ljMY0ci16vNSVJP0sp+s+vNHU
1b5KcTwPamWBsTkZmPC5Sh339Y6MsAdSLL5W8Gfv6bXA7fg2cIpr6q1dQVmyFxN7ULZsTzZxzwL7
X5AUWiJkmmCtm9/reGU0Su5gL9lSLq1NnrYDEKKR8vduz2Jv3TRhrLC9fv1Sy5H6Xkqc9RPcYHQt
9ssdxN5THWxWliEC7fFUo/qaKW9nsMnF3AYApAeMgmDCjMu/9Nw/twxUz4c+skoOvZAOTYuzFRN3
SdRhJ7fPLIiqU9SB66/LDlMPhdxQCQY/gf7BVkt1IzOoOaTR7d41KNfxaVZJMAzGnukut7wsFNWX
cxH8TPDHsgBupk1mQuwGVms+zCsx52Q5ztlf6RwTtx9xs4fUlT/sEAXoQWKICGfXV90+LuEHLbWD
qBELQ8InjgRSKXA16IZZbpt3u3ougiyPkRi9DamXGh4s27gKnOqHg+FXexTVyONh2+JAA4Ec9cba
L1IyQb/2+nJ5TtqXV7SfJ1fqCWvDNhCaKm6i2VKJH2gQVnWSbCfSWF2A0x24vArUiJsNSfONvQS5
gFbvQajFJcqgWiaa/zRAjJ2JGfPYLM4rPOer+6JDSXNdJhp4VkvI5VkhaTYv/MvM9GzdDvXX4SXP
VT3ELm2ETyWhHpEo55NGbOZ5FzloA8dHBj8hgI4rK5N+ZGTqhz9GsuTgNZZoNE9RhJaJHSnGYfUQ
h50EfDw1xos/3i3g/5aEJljhmzSYAwx0rkupqwRuFlt0E2lxYVlf6KyDGiuKI9kGCTWD3/K39HCl
CV/sGc399Xm+Gogoq02m+qHtl1wceeKH9YeTT0BcSDOUcbzTig+hi55q05aNBPENQ3/wTAtdfGbW
xEGuVOnflapt0N+dQU0UDXaUUsBuKEVRk6qoYGUihuWgwGMU0drHJ2aNAWTRZ2V4esRNAwMCO3qg
QKFMQcvnpdZAPn86mpyEe0PVomO3dRiPqvdcBVlzvWj01XlterdkN9SHuEtuvKXUX+ghr6G8DuG1
zYa4Oq9/hXX9YDXLEbXHasbv9lKul0J8NikFqJlxlj/pgzdBy3c5S3DP9YjQ9cqSTVUXN5qi8XfC
ottAIiEby7bTfPkHmhqHTNr1ZRjP3shUIfalaSnHaMuD86RgLQkLzplSBa1H39w7SB5pwapa8hNm
yej16kHyRIF9jhx0ObJOYryF/OFTlKVtdgryTAL8wqTdr2HwubP7Dl7fm1upJQjNMTfCtxaaVNIq
B6nR0swcTYrUsdthK+ZJeN/YdlVGAaQkZD1fBQDhE2QVaKHdQpxB7pTC0T9b294KA8eXP5p291Og
3+aBZaVAnYT7ei/f8pyo5s06aEpyHUQJFTJ430Gpkoyu9GGUiyi9MtQSCbDTgJTFpsMLbla2phma
iC/bpSfAdGQ0qa2/FlYxMp9iCEqEV+OsJPGANcpHDX3PjGkYdFnFEdgbaxGac5Z1BpG7vry7Gmh9
1XXZ5FG698sp0cYsbPPV5jscczlhZvn+MnBXdy/eKQ30UxORuADjrjEyt9iMMPfBL6j8P8YS06f+
x8Qat2/pH3bQoQHJBF6QOpjrQXwRdHjNnj9kc9B0qkGKC7BzNJFxtV6WBM6unoA2zGhLPe91UrPr
jIy1Qa5uLsNZ8v2OU8/R3HTD2eu6ipwRSO8RT2jScALyPMiKcCKmhPLgsiKHbP6heQmMHIniMY1y
HOtHKH4XuCGynI7e8dO+IvIuEOlhhbyMbhC5m6Pdljp/K5P/8PeYhzVBQMO9/xwC7LhncWMd/d0+
DQ4AhVK9kT/ZP/Wol4YBjoCki3EfkYvIKqAj50NthQQpafB1Zu/nziPilQqSuIhErf6n8/p3Yu+M
zgLwgmMDHZJRUwuK0m7F4355e4UNYh7BPOupuncetJ+xmDFn3Ha2pLefCW9x0hETeGM6j9d3gd7z
3AwOzLP2IcxLF/rB8XiBZ43e0TtXAjKLrxwiYUIxmxG+L6/CoI2CB7QBsWhNDVyWiP5OtAz6NnUR
qbxkoL3ujp2Dj9VQRkgTyMKd2/H3ygnGGQ+9ccQil3yYUwiuNen7an0r2EF98swLSqCt59iccisx
5virhU3QACR2SYbCIzxhQr8906yzXRV8/dKzRP7BK+nWN5SUuVv9/a7+uLnbDhSRkMXRnvmUeOqs
G63LOLSiKkuu19Y7YwAbePX67bYlYfQyOWE4lw6ffCKza3Q3c5gYgVBEcTenwckM7+85tZ+Sy5a1
6fHEaOqbS+gUIDAYVNuXKufz/Lz/hGWchMyS/gOYHQAVym34xF+Z021aFA5k5PrtNaU7e1akoZMk
q1bLTw2XexR8tic8oMkfxJ8AYLmQzdz98eQyJmgNGtby7mLQhMjmyG/8/zHJTj4LnWPatowY+Rul
lN7rlc4TMXH++dviy1hSbxufSo4761Wxfyx0d6GphVF/YWaZPNiE2tVYgif8dto+639elvNze67Q
xJiQZ+q1DbFqXKGI2ksZgn0QLtF4YuZALKqirxYrVXAOps5+LZUcZ4QbIa8voemSnNpEqmNxd1LD
tZuNo2HjQCtwnROo5eQgoX3sTss5QT9OAuW8uhz5uAbMoLEfFhbfuRHDh78tzbVtW1HgHI5C6g0T
hmqrTf6Rc+2ycWFm473jed/d9LHPpT4ZDK1CTiI7j7nZ02ye9gwBtlDx5Zw5eEVGpuNiC8NQoDtQ
iLp3q71qARrKHCEPHiK7cdK4SWSaQqBE0LjF0KpXWjBikBbd1gsj5HfJjMqz/0otcrGAY8sYeDVQ
lvbkcE3DHjZh1uE6VsWcRuOwd1jqz+XVfftxKSN78tVVBahGNwdlfEP5ZCohxWK/5k+NPBq5F6LO
rKeTVnrojzpaIhjBBQTAnpBaOmd4Y7VXY3v+q9dlTS1yYzNKN/ecZdIlmkhLtT8YP/WhSXXcncSd
+3eOHvCBOx3zVdzEfifbGZlgrDR+DfxA24KqDsCv9G6onSg2bwxFrWGXs7sJQMxvyPNjASZFzeHX
29YLp5T090ayIgMvtG+xm02lwxf0883ot6eUIKTc+ztXAfNlczd3pEJmnjjIaSUpmb6L+Is6Xso7
n4E436TA7aY7n94ENkQF7yPoQ+nemTkssCrBHNas5BmkeFx+DsURuWOYA0TQilscVj7tQXhTwetQ
WyElpEevynJu/UKL0ScWdR0CmV8PGOb0ykvlenyPq+yDCPnVeeYX1/2yW2WrOu5gp7w7ao3rmI44
jsCcWHQe85VehmcLIhNGUvUbwVHfnKuCIkzMZ/DJ5VkcIMvNsR7y9IgA75ytbtlBHm79GCyO5a8e
UdDtJnKM0qvcBa3KvI+wofqqGZdBat9aH2BJH6ZnlJqiiP0xEX5LyAxgFdwf7/WdFuqO4kHiV/TV
HOVLGX3xmIYn1bxY+w6O/wbPNELURdz3rC+I2gI6MwpqHXFid8AALKeTWFlUIv/y/E7NXW7lvy+k
UlKLou1uc1i5f6K0DzSRDTr1AlJ2TN86U0ENs4YAmOMXflvKhcGqKP0YNFDgsNyW7OXcEcDOlbWC
U0CMLCwaYtHmFlW1p81dMFvl7Cp026DiVao0FtAUiJoMYFYuCD6jdxzifIWuhFuoW4Yp3Tw6zVMc
GaqlvdqDclGXZCoMOsCHCRsXWwwAFXfG4BbGa5eH0+uJldBWrXJBXObv22yWCM7auwflWLgnFw6E
gLLax+SXTmlCPLTBoYbj5kGFSmbeqjqKWRyMblEJOA4wOh0mS9wLTZA4yzrZrSwe7wLteGGl8iE+
WkkAoxBbC6GJok0EjGdtRkiIpy4Ac0bcYRzVKMwwcIWSM7J4ZveTnztyEZPV1rN3mtP4EYFvqHP/
WqzTjVOrhCVgMkenOC+QWKqu+/bsJj6Y7e8owZda6mygPSJ+GImW8W9c0j0kZvJf6SHqw1G0CLLh
OsPmzJOd5UNNg7MXWPe4gipHl8n2e9cxn9ZdrrktN7iRg/7likZyDT1AZmFVPD9/PNidLt+Cv5zV
c7qGYmqdhv4tV1g4xGKk+ZDiTwmISCLOdcko8w/1/qzK7+5nsYshpUqiepN4ZVmOuu2m9DiHGvZ4
v4YC758P+Ykq3odwRiWIXIPoz0Cm3hk29Y1MdT/oX/RIt6+vqBo7kY8rP8Oxb3m2RL737FVVTQjN
DmDFoaVuiKKQslx1emAbOc7c+1Is4u1oAK9WoP4ChwmT6qYAqlaS4Pt7IZEHQZjqCcNtbmK9YMNz
oWQmoXub0znqwubWaSfeysQ/LImtbPXWtWttFkLKQsVvNgArMSM5sT0fA4icUmfUtHkY1a1AHLxM
7NBbs0nHpt0HDogSClzTRF4IOCENR5pzDQxAHR7i2Ebj3RXvBPNXz/M/RdWp7IkWVp6wuNikZSo7
27rajl3dYf0rFt3EfPfyRcnlPoG5YRIuXNdQmm/oyjP2V8AmmHeo5/xp1+Fy7/9jc8XeGRAgQPrf
iiqQGgTlG0Dp3dsfxwqhWTSBt04Tt1vFkcZT2rcf0NENkpRHfr7BvhXlsK6KmkXE6QymMZpaSkMM
0llH03Bbn5u5VMhydLUztIBMsjxrrGmbRmCL+tLeD/Hj1HOhlcyeO8bZR28SL8y2TrWOCBYCh0Cr
T4kT4xRJ4I2IAQ3D7DyJLxZroT2FNi+jYNKHRRlmbdGlQJmoN0NJ/3QYdavsJKiAN0c1SWn8PzR3
uplrNvVTkVzSatvfKY8CHBmni5BD7B9mLHinYb2axdyPne5ns3YFWgvm2AW8eu69HXn6qqv5PaLq
4YwoiEYr4mj8kWYJ27fT0dRrtxHnLzgD7Tgrk+WiyuU//RgFDR1uBXL+IZHp+YErR23jEWuzsn0T
VgfAwjNWt+SmHs3T6ZMItlsnSAugeRcE7wxtRcYGo17qUKKENEO7OnMZpDcFstMmc2WcKJjktXCQ
2Sr520ZmJ8vZOVQydyjETsxdsGGYNZ39qZXDqAZhqQg+zHR2kvi8IhzKy49jMza6vT2qsQzHBmSl
fir54GEMOvIYktkoDhiAMd4p3N2mvFA6zO6QaktVsFGcEJBADQiMWAu32JUGDnSZbORyNsE2QzvP
GQgjz87AYg9QTzByMdJvTF8lAe7QqUJHL3AnosY6rYY05TmBXxMlT+vZccoOpHwR+YlCL2Q5IM6A
lm6CQydtl0Ep6nmzxjX906e5Kf+Ypva19NPYnPVcGBMr2xgqmvog4MfQjyQ9ZQ3B/6siCvfsLslY
l1Njm6NS4bV8DAOuiT+B69FFu7FJtEgY+hoWi/LDzIWwHaO2ZwMl+GmQlt0wWVEH1YlMu+t3uc2h
Zr97Wykk4VPpz+b0zYbek6E1uz4/U+QVDy7xx8C2yiIhjJHPhZ0RAzRlQe0yhWqJUXooCzznlTY+
PFiAox7xSD2s31LwBWu3uNPFrLSYnL0kkDlC04M/7znkNaLyu27U8oYIJKYsVSZ8e3i/mzIc6VL7
vFT7Dpfy2GwevVFH9dkU6hKF7TsGStTy86wN/AtVmKuHSqpUOfR8B/3gByet5aiFLkqRoQf7AcCH
wn0t8kokRKvjs7CoVD41x6EyvFF0x641qM26iQY3kMxod3ftWY6ZGw6T46YJHA6oArY3BjpAudzB
rcAn1cqH7zUmpERL+Y/oYQO6FhGXIz5xpfDOlcAhITegqYJr8xTIwTizKMW9aGFiTgLOJ/5QiOiL
iaMqaal86q6YZkjhJeaJ4Yxk0s478KAqErB6AyXjRC5VxpN8ttoZvhK8A4HMVtFE5ZicFHW+ZNUl
M2/lq8WtZ7C/juI54A8ivVV+1aalYGxaCvUDIFHIQuKhXTxjZMHvjlVjkqvniZCMW+jQ86dnk0WI
EKmBr0syP62YzpZ5PUON6D92VgwombRSWUKr8v70jWzVb8sA8rTTQOkyw+W+UCklbFFS7xHeyRNl
NlY5TOuUIokCw8TzOo/XHrGlNxe95wK7uAXLN1mmojM6x2oFdaFowbtF+pCHveScNKB17XLDsVpU
9/AXWjapTFFhoIEGJJL+wRyzd707kI470WUfO+4UJhXXXGerdPknxr84bRFnDG71nl/7v/mfUPAl
mFqCk3qC2f+gI3M0TJyj/K5r0FpILWuzaryUirDxc4mRh1KalRs4At9r75paUww/MXosos0WFlhL
rKdrAfEBKPN5Ro0XFZdFAJlGuV2Mfk2+361WRz8GI4qxhP/rwT2P/ahsYiJiCHdHht6q23EZUHIV
38t+SX8YiC3sdDwozr2M68EtAHi8F0dax4gHwTIQhvYmYoMUXJTzKevcOJAIs1d2nY8AIeZESfrm
4MOHLqmC9kyHIUJTeGyeYEpbB5xfnf7v+nBxPWbLGlZEy7QxvoFz9QEyk9z7GLotOmU7E3vhh7kG
bQt7B/BRg9/xUu/nRkN80DsjXhhWmUjpbfPEQu+bOs6mIyuXhhwa+ysbuwtEHjeEzQOt8qK2xJ4q
SvDXaaGtVJzKe3Gn2v0DuJpD7dXhyBjGlYTz8iJqvXrHt36ofkg3FCkso8ONhALEruSy3XrjvV+C
zHs0MOB0SdM5SmWl/Eavs6IHOWVM9a/durDvyn572/AWHbVL/8sYhTSzjT89yKeogh+DMgMdknDF
Ys9NQ4lpyzhs/J8ooVnJ+hneYIpGcGwFjp4Yj0Ubdq0unHGocpbLdOGLRrFa5kxrIfdhHbJdyNn1
8biAr2cNJB1hPqFaNcymqWCS3a6clfJMHZG07EoMX6p/vFd9B9a3jSJdF1Zas+Wk0M9tjQHEKlLX
TAnVuJ1W7lyYjpq5k5xIjcZA4J636/1RWidPqFYAZ8oBepNOHk3vZvozBefHnIMcxyOoyG1QQ4je
djLoejI6TBCovqiDrcuWs4WGgYAsPvDUMmsU7N6fRX+SIrNsYh3LMtwtRQsji/CmzzKR41o0TNth
6wWV9KnYo17ADmXnAVYpfUq0F98MIzzsGsHbc67pHx1dFoqOhrsXzRQMb2M6IM/eQfDUhD3IQMlV
wE5NQW9BSeI7W/GQqGvTFBFMzGOt59mtLOnb7z/isHb3nxVmiiTB810U1YHV7m7ZvIRJwhMwcWjx
xN9Ph7npQB+J3PmIQ46v7qMwFTH+T4yYMXH+cVfyIGPXPgXHY2u2vjC3NzjEH6iPmt9Bt9Xy138y
Cl5RImJERGvFTmrEoxsOwiOOpFazWpDWr8qpEx09/5ebqp/K9hcu09JRbNPtayF+lU/hsSiajUiq
K1WdLnH9lEAARw1IXyhHtQU+aM0ebHIRcPWq519hoaKklkDiuMjRG1xDmNvqAc7Ekm1GKa9lhwHP
xpzYl/PtQtqEj4kOggdDLhNjgHjPyj28494v87e6DbXAj4071Wf98GQ7mhe9DhNwrJAC9gy5d8wf
YXSmehrKDrxcZ8x4RKhvTA0hzBBNdJuSUvEAa+yBGaIfcyyoFXADS4L56q7zfoao1jnGGTuSZ6h7
yxjVMF9FMh6jiUfsUuiS+0UrISJUmor7y6BFa9w1hAPUnHRG6ItI1TYuJn0cwi+T+ne24xik7kkz
nndOezvYQxyF1bmC8gyt22F2OOfmoOUZsFsjUO+qZeI2l3h5NNSG+iSN2auBmWDnD0K8aXZkzuru
gquK5ZCqijwIqLPTQS2jhUEQeHxajpiPUlw87Xaen2nbJJuJAG+KryS8J4D7gBFE81K1BoMhEO7T
XML30Zal83VGlVuP1MT7QiGseEFBs0y1JgIZAuyM4CH5f3d9bthepQcd1flfehtHmY/m8OVR7N/m
LpZnIvGZjI8ncnosASoFUeteRmDo31qUlR/gFXO4uqTeyXNhBjwE2+lz3LeP4c8yN/xA6N3T3r4C
wUrWy+o/nFvW4GGTuDf+WlwRYqpM+Jp0dUgrW4+QqryzYPtwW1fPBG66HNIWHhMqIj0FgwMeM9L0
Xz+UJGL3HTA+6vtt5/hbu0B/IL5V0rdJpDDjIpzszV6fwVvHHX+Uby+9Sf4zQzUWxvL1SLVuumGR
RAowmTJSijWpE/e3HmNkO1GzF2CBNeej4Lg29seDyDBEkoL6/Kva7xC/x1zg6lXkwF2dtY3MCyeo
diAk2PLbEi/Q9XGAYvKKKll04iLwqKpNW88YyvmbAwg4Tm+9MmRcgznN/4MgLv3cWAcPZp4tml0g
9WdpV/6XcBuGB6kh7DfvhyvJJ+JF9o4RUPogRljOiM+ea2CMD2sCLTV6BTx/7J7120voMLSkP/Zi
jleFyED5VzyisF+6i9qSWqkAlCDQI97On1yfV07X58LZYV0/wRetJwUoHgZ26+RCgKzNMicmtUpX
Iv2ChQ7+OKg6db0M77z5yE2AP88fwvix98E2p//PvwDqHNrF+7YNKjbQscyPgH/jSYoCz0ibK7gI
HqxaoBktOWRXmKl1PHa9kl534ZYeA1PoRyDDEn9GOon9GOPNW276Bo8wtaYiwCxDX8ZWuk9dyXD2
jJLzVzDiQ5XhaNjGzAOZ/LEW2Fp0YvZ1vjUEbX9jiT4mxWKl5xS0tAQvOWjgQcdb7Jgroa50zpa2
gyRA4Wu0jx2LkPTjFTqASQd3FsKJoBXTWujzoRZ2eoIIsRC9/RPu1upltseRr0SeHjjFYxFsZ8LF
g8cly6n6iHbELi2fmHvsj80OBnBfPCJNTaEHf2eZv5EmuvStHnXxwkwzzllk3vVl5dHPXP77UPkg
phVFsY5L1DmQ9rgW8pidCDupYxaDB7y/5h6S5LDXr/f3bPDrvmUVlahx3Wd5X2gJ209IWuRgITue
+x7+a/CktL8tXCarTOYzjjIiA24MDEx2lyhYnf2nLQBTLRF9bhn84sKiwnU/5+t38503AvM4asQ6
tRRXgGWieyYkGjBJtaVLMjpXPiZUx34Ar3/aev6SIIt0bqsQUsOd/e5edgd7ha20eTbOVPDgPynr
9v9RPAryrUUy23U84uqM9W9NV0YV9LYw+WAA2bT85cLkzuUhne7pW5KvDxI0WQB1IYZ6zfJYVEZ8
GdSVAcuhim+y3b2oqvhowlmbM0ypJ1jOOP+CiVjfFKsvxLZZ+sPVKqdmmzBe0ZaVJRy2bqS8Fvpy
3b6pHGJWpq7VglQ6ZqAJuTF0iKF68NJABA5FG7z6NGhBZQpoVJ4e9R9K9iaV2H2Myl84TLw5w7yo
MleZmtWkhX9hE5lQP0Gmecc0qcR7v+A8BrCa7ibVq0p9nCu2GHmtRdPUll6xU8VV+s/l4A7IDbqF
KkCIXwDKJ4TTEtV4tGpAyGBBgAwKoN5ZRZ2VfuDJ9Cc5tQ5Edzw1d8UrKbSx7mQQkwW7K329j8BB
/ES+BUg9AQPIDrmhcic+Fk3shQX0q+ktFDGTGjsYG8F8SNtImtU/rJUU8QH2kBoIWEo+MuzJEHmH
4TFrdbbhUzxZ8FbhoOqr9hn4K7OOCiCUhbTGXOUu1cwXbKXsxLFBaK3o1Hr9/hq72v/k6GwMuyWT
w9kplh07qMWdz5asYwAsayu6KdOfBg61TRr+8wNR8vmOLc3T5v6+1x4dREGs/Oz3MiBW2L9/AXjQ
hsBtvKBPt4P+7GpXxJahyKTrr657qrSFtP41vy9Xli6uGrhYgwrf5bgDnUI8Tdi2xaq5l84TG7Fs
9jpZb8DKy0l2X9PKfFdr5/RcwtpcDK1vsZROFewva9b/lZ7iUXpNeue8LhYCryu60aGMAroNxt+o
xUYbVjRp3rpM4suf8uUg/fFf9pZAh32L7kE07lFrRS/zztFhHv0/Z5zJtyVEDr2ok0MwSVmCtbzb
yMooRzHgZDo5FhnQkn4cyC2v021dhX3u4RB/83tC3Y920awgT8YvB0XPGW8CGeOqB30yB3diKIJG
r3qu80JwhiMgUnfU2adbQCYQfReNZdkgpuI1y8ju4rOjtMpF5b1xFdTUDgSyPu1kYpQ6xDldsOjS
9YUFA1WhmezTWopfKvEbRZTRxNOgrnEYwo7khxvRLHcboB5SboTRBdwQ5HsXJGPdtcF0+GeloyrD
fPdU3gLWhOWJiP6udeNtWgOy82bCr0FKbYNNHynI3U5KdzyLvS0M0OKrEKpuWgdqQ8nhUAVj8gLt
y6ke4n/QD3vLZJUz+XuusAscqtq5e3OQ4FcHzPzDEu0WUcgoKPDfGv/zdSbi6CdAL7x9FgnE1Vr6
KuVL0e7W5i8kw/gwEhoQcqWgO1hx30bjRQxvJQdTu4FUTV+bFaHMaOfbgzoShK9e2qlRJTcCamgQ
n4oPb834GrNaiNtLE0gC9R6z7McTCsagHc9Tfsj+1yEw+8AeuxbMZCOTwczpVNznvhd5WyE9TeOU
lqXh347RA+rTN5yR/t3/NvaiGZGQ98QOExsMTmR1UreS7ocyL3/kv3kc5lTFS+fnmavvm7hZLLCx
0ioXdCRZtvO8BnG8u9mHSgOrELozii/P+74w4kwhPSnYX1hI62WPaZhbluddjZzdVQBVIQOoN7He
4zVc9cdNpfmxPYS5s1Stfr1zQ3HMhDk3SkHsbyiFT5w5nN/RdGDkOU8T7g1f8xix9TTkjXi5+4al
wiPdmSJjEYvIwawI5nGrAprdPVoDqma90tkbXR/jIbLELA8+gt8U/zBVOgpKym3dtHxTKGrDTLvn
49EWylTlZZzsKY8LZZrVs6164lfIWWGWZMKHFovNWFHkKxFu14sqZOJut01aZPsyarSvtLfsBSSn
rmIKN8FQOmWzm0pTV1j59YWw58/r9OMjXnKn86Wz118XvCGJjpB7MqbCqiYv1HLd3curdwR0R2VY
i+KYXolEOBXmXOVCcGkDMhEtPavCbzYEyvBdNTUmeLcUw45YMtOhnJk0KoF/rM5ZGUdqyWGSCIUJ
UCIkg2wfK1F7HlYH98rVGzaL9xDB4HyAlv2+ceUeyNbKnZKqfiBKOHbmwDfkXES+gxf1b79Gf5QE
52zlUhbLG9vD7PSazTAOe8V5WEwkDNy7NaBxvoPBrpQSgimx1bghGJ8x/xqTdQ4JdE59BGQaT+kD
CVGBzSGDlkIIdyiMyw1PncPHYKzll1V2YIuzu7doDxqq5UYx1XsPsB7m2AKL46yHTZdgEMpU+WlG
FFYMmUjM9cX5kYRL6NJUIfjyv45E4XUsNXEwQe+oekGDjUOXLNdn2QpAaGpsmiNtonp82UVesnen
zAgyvmPNMfg7Ds/cO7qbikchY4AjhL3hKtMnP3r5CKqDbND1Gd3QBpJeCjJ6sdnlLcPgR2HaTsHN
0Y5uMLL8tQsG/rZodjs8Pf9ZcoLPP9cLHmyXnlU26K7iYf0tZhFcHlG7li3JsYCtigCyHz9uLxbX
s3f/SVT2llmyD8K3sqB+oipkzP7TChePIlXVQSCcrHjs1LzEAPkMeO0tzucrMHmHCAv6m8RMUUVA
c+ejXA7HDrBFy8pg2xtREUrg22fVnKVXSWlmoGmQ1zD/G+bUVMQ7xXiN32dhfxatrqh+q9Ha//TL
hcWQJLfX1/Jby1DMitzIpICGOEQFhZ0CMMa1OAy1YN1E7j96PDqMs7f/v2EgXNCJnPsP3Pp2n4ib
d0UVXA5mFZ89i3bedszf6e82ArFucpzgHlFE+a/1iVWE552t/6pEvqBH3eU7JtfP4V73rJA1I07Q
AQBV0GfUMzdDvr/B+jvioE2UhRYPpB4TBK8M5O9f+vJ7stfTpCt1VDD76OBm3mxhbfDMAAm82ufJ
bxD/eJen9XIg8Ud1I6eF2iLujEwIAXc4TOAtrFW1bZ5q9X8KhBir+43DFEMIWegwbZ6fzq6noD5B
jeSs4x4/MeK5E4/bn+txPUsSSocPQsCtk1KXiuXLlB9dEu9zgaacuEgbVi6rs1hw9qrVNqbfPxvc
/3D6RRYmOCcJaUCeagMEr/C/dLUW6SzXV8gROCt2QHivPSmymxE25rgIDQzByVQAv5ZIR83Hh6b5
u1++WN0dYzHwaCjAq0a/EUeflWPFvjq/eMNwRewPEFj1pj3OT9CY93xy4ucVD9kuB1WwzaxP1yEk
dk7TBCaSQ8Ldm/qrw170VnDdDg3D0cIQJoXG/m6BT2FQ8unn4r+gLLzZ9TOIjxS9ax5u/WGzAbOk
Y++Trmkjnt40dDRLCHBiBBNc0PJ+hx74dfDpreBvDkkN7fpDvG+OIqeJcCZNH7lGmwVPp+UykiTF
xhqfA1cTcma6D9R/c/v1n9y2xWKtxZU7NAmrFZ7uyS6Z3CbXYMX7+dkPQPhcnMyryLtsZvg0cy0r
rV2+ByRrx9RUsAC5M7QMf5pl65Cg11U8uKP1j9gWjroQhkdKi3F+pM8h2X2pQiagfvwXV7nVccCQ
3xVlqM9vdJPa/3yePlvL+VBfnbX3Z9H7CjQS8z/Li063rgQ+SSffOKZpchJZPhCZut0E/2rq1qj+
DUPW2z+i0ey1jdTko1UH+ys6IP1ZsTFYoDxkOG4qkgu+TEKCvDxem0ysm6Ue2BN5/cgFa9KPBb9z
zPECza24ueWFeLfAEMWBb0lkzIaRPp8/i5k36/WYoZ8bDDA9w8WKdNkvMxSKoeF3OZLLvvPhqXqh
0ObQE3WNOy8aQniib2Vujf6M4CA8TB4II6B7yLJJRYpw79cwexwdX7dB2tceClyqyNyNCenEIDUt
H1H1a+JlVGHwxhCXKDjvu71cctEzhwsj07stwxHcaapeOUWAqMYs+SxMqSNKci6t07qJ/o8OlFsy
Gv0rgHpjLI9Ad1DS4EYOboJY4Z9bMlVpTgPQO2RIbYF6Wz3oUldfbljXRzcuSYli//aGcDezVkb5
E5gDlyhIluo6YmEyFSVm/klJmgQZUDX10BTLDYz7c8rxBThxPAdaUe90ti3Bi7sVhc+OP8w4NBWs
pLMR/FfH1OCErSVIpxgVrQTveFfi5oC/Wu1Xb+qqG/EIKsqviqW6uT+RFfoctyfLY2HsMdzknr5w
n9tFaGWrnnh+QQAX+6eUmEDVc4+/+V+56i+Zp07r6xKrKmLIcubtndan2en06LHipQE6Pd/kgq/v
v2vHC5NWDmCfNLE+xxLF5cTcK0Oeuxn9QxvRxEJkIEM0Xqa9/EU6Zl8f+Zl9vTjcVnwUAFjikQLm
TSQcZn5urO3jbYR4AM+HRnx91Y7hHS0veYqVG6x6kgbWAxFCwwleM8MQbrBB5o5Ixv8Uqu2Sgdu9
pHS4d2Wj3eUISimc5EgA8S+8WBLiS62zPX7Ek6Exf2p/gClKQl5mnnS2my9aFDYPP3qeZWO+8BwY
niAFCg4LzzzqgDxwGiVz0pgxrvt98zq6IhCRHLk+KzUgtRnztyrNx7OypVnQRULru4zHyn0W3h46
IMj0ZKe0L3dveWdbUq3+yiDyxZLyoe2YDbEl/+Ca/Nuvkyhl9XRz30n3oLck53jMutNFPeFpiHBh
5leUbd7HEfZO7I4Ej/k9qcSH8aePmFEFl2BjRo/a2TP41Jo+u2gGjPuBo4MnGF9nVA+sP8ArbvNT
bO+33X/FIUfYu7TSQepKljlTMc4fYu9uXPRkN/slRMqj6hzoTF5ySTwXQbUu5/NhPAUZCNMiyTVO
apHEQuAu9FTVqiHbPMRWWCJLB3RP+eQKf+0g09kTPl5n/eC64w7lDfYt+ORuWktp8GJy4Qg7ktIz
0Fu08Yqdz9QQ7w1uk+SM5mgGWjR/0myKG+gn1yakWqbsIS0C/u83OHYmPsdlGWgzqsn+031nl3eV
33MuCV8C0BhfOrYhMKEN481odgJOMpfaNxEKCWOVAxVIMK2eXacMJMzmdUDmJ7vn7LN/mtHChKIR
+s7K5ctwRFtygd6Vv+FcECOGihExPscU8beKYS6MEO2C3E5VRO7tEDx810eZ5hibE2DIBIBp1VRX
VQ5bVTXNP5Mizb/Rv5EN+qIy/wQfr+H8vNeKLtbkShoU3v0F6Sr5MsR1trQB1YxtBt8+oe4YoZ3L
BsFzs28UnhidlYbTfOFVyC9DtlQZ3usWswIqBLA8XHOrg0uEhxo7I+IkGO9wj4u/9xf03Gvjzumb
boD4eZcXbhh3F0e1nqJ4xOMVsmmXS3so2jOGn6SfmPXIkj25YIFSia4EcIzAmkbTFP1l0A1LN3au
YL6nQxAsljjyi4vBulwJn3HxDzCLBhwO7DEtRlDqIWX9vepkDeOLctqD4VVVqh3zkkLqFFPwHmH9
bzOOq63+4p65++D7PsjrE4QqjvuFpbkOWGEcohl7OMGX/aZqICSsXsnY1E8hnzW/HjswRWzkNxus
fqXVTcESabGDxHItBTJ2lb1qChMXI7YzP36SOkxfad6cCA5w6At6LP3ftK2/P1tk/cwC4XkKuPIa
+klJ/1q6DiQI2CVdhwIvx3ucl3o+XkumpBfKrDAvQTLCVsV50Z1LrO9cdSVcTHkkUmBloIqwhMGU
gh4IawLjaufMBxpHqjnz9vDx5PFjliJaiTOi23Ks0AmtLwCbTVO9DUEVEOFkadpwWwwHeOmoSEVC
ivxF5JMaebkWIekQKnmqB/bfwaipTWlcZkJ4eTVH3zOuceCJTlZW0NimzmttMma+ELmvFi3Vt70g
KMl/1IRG/WWl0texQ5ilvUowEttgm8fKhHRSiXNmMiw5j1GU4kigby/ZG8+ZiMuymVLmvto2IVUJ
PW46+yp+eRmAo5fUObaV6Z+bxkhiOzHKYN2zQUvCjFQbVSVqbBX3YPE2QOa41J4Jj7j8d9OlJUrX
ozPxSw/XZZMDalikNV7JwywG/CBOw4mJBeWA21SGlXu9ysUlKd1Dgrbahaa2rdwSgS9VXk3h+xhJ
dKdvpyysmMtmGMLM0RU5lGPSsRFUCkvIMFnrF7RC6njkaPjDECAA48zyF02nGZp7vyrlmzF9Xyxd
mLEL7ITZT/kEuzkyvnnNZBh5sEiD+lfMakZrvVHv+SxnehY0N1wCVZOLJSBqUordGdqopE+kNXil
xFcyzhbvTWEaCPEtPd750oikq7WDHtoajbedx1VFj34GFOBMOoVjL7rGy7R7Z9YSEHFEbY6aHabW
xFSzJr4o005x8DrnnQf6WaRa/FUQIcHZSa9n7RnAJvIpXqPOjfPKpI7EawGwsUEbabnolnFlrFWy
6AiWYlVgbVbyqkA0kRPJQjf7NwfEbk0JrP7b7rrYRRwLqHbFW49JkXBBHRFHx0vOp9HkGrLKNgMG
pf0Ur+HjdCOnQi34gqUdbiEwPyOwhe72ACfDY9IkhJPXY5OwPKl0b0MDaCfrZj8OshrlERYU1Xff
MdGA2kAMNm2c8YqKe8wtHXmJLDKWTkEndtMLjPl5nM0TJIK9owpLrOWl7qKebvVZ4mNVFkpwop75
45SdbnRZ1Kxcw0Ue6BoJSioo8oNdyFVxy+iPa9zWzLvmMlWpAKhhFIqA86H7G5RSHbKzrmTqHtSU
F5jTH/6yMvcqApMrSPzKokz6s9RQs5KDmA8Z4lmdZzk5nX8q4Hx+6jsyshiZjch8WEmyK5URHlnF
lqoRRqnrSTsOZtn1Lg8Fzs72VpHG9cFebGo20v4PJeqFRJYWgdJRlJcKANFrJUnyIi3/K5ov5+Ez
KUJzwWgIPXqGw8sg9dfwE8tggrsTVgFObegD4tchaPkVMKWeJMz8ErXun0c3Ja65vI/ftuEjwOT8
BYOlnIWCCkqnmjw+n8uz7awtvW1EY9JqQjmGHdyPTRgLjTg8jiJueT48m8ba3iU8dKr4/P+I5hta
ZKyZQyvMEgema3yL0gUCj/EzOY+jda3duC46wFiTxK8ahlCorvf38hoFVdTI41KB2fvqxwSyixia
oZ41675kDQAKvnsp9nxn8xQs7o0KXAGcAT9yvTkqITYXcDFOf4uE9h8JMgGJS8hpFplLJvVXbxOM
i4nkMZ6lB8m8PqSrcM3dTNdp157lsvSwyXV3QRAtdEyiqgZefbcbfqnqXMNdQEAvyC4ziwX/mOaL
KKrZ3ozVpSfQbCXbXJsBp3S2zJ8BjCTi2YpTHOdtf+b+HrWbEpejH7+cXv9oQ2yfA6qkVPvsUamk
b3fdUC+nk/1CkWbFSuYqSj/l/rACKvqxg/sI+29/jVp7OLWON+ba/PSTe/xaI41T5MRYTmqKq6LH
FAmh9+HM51M8eALJldAAoAKwwDaVJ95SlcgwtNJ2WfNaE8NuiZL99ZsnsxktRM9PINQprivvFhCI
niJAUhpC8qR+PYOmUFrcCnS66TrDrA8VNJY1uSiMeH97AUNz0pBBVdVlppsXBjI6vazYZxowX+Ve
UPQHis3ojyOGwkIkVdvx71OCl3UCa4CH/zEXRuxRPdY/Jzb2uvttl1MIArUMpHhaXKyUoLCgDsaj
lVSG7MdCjd4j5joWqKTMaYNoRLbDJnDG7dQn/Uzhvh6yjSENtmyWLTIUasNFat+SJLTdrJq4oNk1
gqQ241RpngLKNKM9JMdmHZErPrviecf7oafA6IPNrVjtzpaJLt2w8DOmyfVd1QzZdhumw15oFBpI
pbkyNC3+5j/47IYQq1amsy76RYoQkfKIrBcbXDTwoe+e6pSVd2ptJDhApmxg+6mi+4bxa/myb6Sl
JVHDfgNFhrM5P0LHaG9hE/w2mwuBxnH2koQREbcQBGfItP6xxVuvyAfI/d0ISfdy2hzkadTAbolR
dR+tEKNYZ5oZUUtXaez2wEQaCaFR8fPT68CmxPP/SD27CdkfWGNLXbdLDKU5noZIFf0/c+gdmGRS
T81jsJWp348T69yjwkztRU7+utfoJNHSqs5Ahsp89DSUED6QsxWdEK5FCMT8lgIrN8TTDi52+UV6
wsirU5QqH8vWRIJNsky0zohR/0jxpOiXWmant9AQpgWWrbeeHvOL3pIIDqO5172vWlzzcbK62lv4
XGqM1sewjwXigTfZak1uAA8pwyqAp5Vdw8GRT/OuiiW3GUKJP5mPuil86BNEzF6GO7fQMGxxG0d4
vOyPAMpbKkIZyExrf+F7BQNFbn0i1XIbhWsNd1j//IugCilf416RBl6Qu88KBKP7IaOKlb1Qps0i
TEokjYMN6u7Eh3TJKABcjNwAt8PgkplsICYAj9l006GURIBHzVK9F1a9jnUMoUrjXYd7N7by9AJf
XWwgwolbNDWJzxPr6jJJ2uqc6cFDDIdn3WfMIu1MDOOqZeko+sz9d1yt9oUb3OvEzXEmdYo9pGyk
m46ZJaNOQlMSnBD7AbGiilecrHk2Xaqq3DMuqvJZ6XEx3Ad8opNCznGc9hsQChZrT8lqAikBoiE5
eHgATet+SW5EZYpIfJqmMSJeI+u8vV+ZkK4dd7tH+uk1wRc2id4SdQsLpENzyC2gMdZo397p2TPi
imn7NCXCQ0KEtbQkoieoLaSNWQZVyne3Q2OZOMwfTOFAz96PGKt7BohAL4DZSd0MV97+JPdfvkd0
qWPQjWA2th/RcRgFcgb8ynJt+DLciTUSU6UqEIwU1KreMaFg7icObsUAl+9uREXhlVIuYAZBxl2R
jJ0ACVLkpKtI/PZdd4rmeL+vDqwocCOwhhZgx76clxnMVtNZsIlPAsLVeV2Gk7iBoCfAfA674Fxv
CAFCL7zlc0w52njwr9SlsC42x1jSLfbNWj5cD/Fwl0hgoFAm6aSkqj2XukQjiqNVhA5k1DBS2ZNY
/1Nf0sViVS7fxvHKUI7Gz+WLJGSJgNdYKP7HklBc780OEAeF1JkQUDWEl+q4LR6E7WijI5+EDqd2
n8Q5waNnu4fDyOdL7VSh8mbqDHCv8N0d+D/285ah9zTailsoC/bTNc2Ae7iP4zqftz4iwZJTfgDA
blnuMujmultzALLYDXup9eUjK6MxJw0twbV26gdE3YKXnbda8eK1NT6a0IiJr0tL+Z/HV218ZKg9
fSjw9fwKDZuuCP/IT6AdYwI7ZDek1uR9TteO5p9DvPb1HM+XcjQ+DLVdi72ufRutXuY1vazgmWHv
H94QmI7+U1YzrN4+oJzc91BbaLOWNqdKTP3zds5+GMyLPRdnIbuoaj5FVrd8jsFcvktQ81rviti0
1rR/hbSuakLLZi7/hggUbJv1PAia1mcABrrNnaQ6+GO5Je0hR4PlrfBdoiYrsL2jOjoVzsnaihY6
DWI3aCZq86qXyVYK/BHBGTFmH8gANH6PLTrbzxA6SV1yZYVzFALRnAmC6i+d6ceHkiJ/FC/CxSOt
j+inLu8COW0yT6INlGshlg7MG0kpVoIAtu8JBaWLkDzJHKdAa3cMThBFpT/+d4w1uywj/zVM/C57
MXFSlhUhoGwMZQ/nvVS8CisODDW9KfwSwoZhvcrCnKOVfEx7N+UGUnFPgauOR1Rc0kBf/2cNINZ4
084JwrEqhPQWHICxF9V/xRzKHhpD845cZpAR1tM66qveanHLhH+78mBZR1UF3TZooUHX3oeFFF0G
aCdlrqb8KfClsb88dYoftPrlBfM/qnhGljz3p391hrSaCjxw/dRvQ+uTudjyKrQaPzU6/mODtmED
owgr40FuMn8bYl3P10Fzj9R9zTmzN5A+T98ojccchTV+cd7kTDyNBfj3dXRyv9eJp47bs+24GfrR
Lgjo2jwPtu7JuuQ7RtL+GPo8hupTa65Mg0UPbAXKbQZFPtsh3bwkVeX2zzv5/Ln6MvbuUhTx9S5G
jB/IXBHCrXUsts84YRlrKLrpoM7wfQ6QmQERvJtqjw5LluNnGDQkPc6pgcSQWEF4VdjMfQbwWwwH
4/5fiGhg+KF4m3fyw4k2ZWXeUQmlgRODFcRT/Ugo21k/wmcNSCLCJjiMMO7Yidew/6kNnELuBVRf
uJ+MIdnzSmJv4k2kQiedJ9xMGqwtmoGZDvj7cvWJ1kixLrnqVWFjzjGT8ES17bQDZpFucYidzJox
7COVIBphak3BTxbCb9v54FIbXsUmJRi8wndxSz4pCyv36DEWhqwfXE41zkZcsOmVRVvSVyBn2d5z
eUe++836atAN2Fi0rZ0WD36ytXfoAHqFXnWlyWIkHLZrVNsdbIFI7lm37nGcdonQ9eDgv1g6k4+z
N1Y90DlqA89A3+EFwg+G44DGsuUvUNzI+K1+vGs/fraZhS8G9PfVuAGgvgTdnL6mUWBv8fFId4Ih
Y0A6Yyh5BuSuiC9vWHTvxI8WYsjdqZxfyV09mLDJLL2sRDSrlNPHxzmTAce964NpER3E1FzXeCRX
GQymfENZDVw4QD9SJT12+NHIzg7/mffKGxLzO7sxO69JcNPov9s+6aN0kVpOnnIrq6vUyzZjPR7N
PnWpHdvKEi3KJXTPHT+DuIub1zX5g06wHb7Bjlk6wrEEYJDdEC1lsHZW/8S3Z8DFC/YHFNXc/tEl
zeL8P3MUodfQZoc9eCU40x5h4T4FolvukG4CdPUxpT05XPgAcHIwkepwRdNrT8tlZi/FDGc8LKz9
i+ttyaP71Q3Q33eSvTECGApfeHYkhxb8FQCh2gWGLudVCxVl4LCZBmNCCrkamo+3t9YKUkxwk031
Flujg3QEAfpBAq6KlaWAd8f7SHX3E4MSohlkTblO0g5aGElJiKbkNmVe7DLHgwb52eTPDLHy/PMm
WDVJY+rfpMRfW1Z6fb42UNspVFrKBYX+2CBquC/52HRK940hVj8+5R8zvJoP3rbtqjClwHOq5OHR
JoCceVFxwpUAG9F9BSj3LcNGbvpkvfAOiPaw8Io9kUgL9IsMqJNMhC/LFtvE/luoCI6VFOpoOUpP
P5/WYQXhMIXzy++KmDr+h1MbnPwrePqVbXlyTfXtcryqA7pewU+C7+iut8ImTmZFE6PD92Txjh9g
TKpo/qPs4WLRnKrXNDFgVjtFCuNRW813PUew88SISivG16s9WgdahSvGOK/8S4UVW2l6xcxxk0I5
BOE24wcBmMYlnIhc3pniL7n/PsjSJijGwptMhB0NafKj4JpTO5t2LcCYtrUi44lXqxDkptm0g686
fBy7HFLbSYOBP8dx2bpHW25VIuioTUGSgExI+RscQXLNznEgOhkBRVxO+KMrugnjXfKEArOnxRWZ
gFl5s94qCWMvqy77PTCfm8Rf3WfKw55migdvWW8tt2Q8289TGwC7CSSPxMiyHVX3Q/5Vzbs8I2SU
Bk+C3fKoqBBr5FLcZJXRvsPNBh3kHu78fWVWGc/7EgU0/lzwKq5leMKc+8T6n8Gc9V1RaMzp7wnQ
m1bs0c/MRcN8ZlHGhMtdvkRcDhGdJi0/+wFljK7H6mb1CfPtyJ3BZcbqkUE+k16vQgJBOMGDGSYS
mzktSCTKrRqn50ezRGKuydArP710yOOkpjR79TIg+3Zm0ubY/16q/Oll/SHwwMaoA52i1SoP+rQP
S4YBtj8o0U+HoU6pX5L7dnRNcgxNCKIsqHUsEKO576TiKlPACWxRv8hcOCd8xhlejyGuyt7EyovR
wM6IvpujhsLS/2hCca8AmP1FrPeGRAaHSZRTYsqz4M75/taBc+o7tGcb8c5qiDOeZE4yMti3iM6F
L9vMSU6e5IHMvCaiT66lR55Gqtimsbc3GE8LoWGbYKtR5zOiNynjRqh5319NZp59v/DEP8KeJeR6
ndsZaTZRZcY6kXZ2s8vFgl8Cr1cYFEhKd8vWN/ILmKy34dPMd0EpPn9JjojARdBv7omP1Bi+8drW
K9SiSIMqeoARb2ieq4oADXaRF4u4e7l6oXIwCDaMbEcLVm9r6ulMUDvvzLBkLV0zGxAduLMlOoO3
LADizzTcb4AD1kNuoxD0yKi1fK7NAv3IJWPLybKsXvlMAwxdbTNBhUoCUi12WqWvsdECSHLGr57/
yrz6B5aafsNKtKNnzfgntSvAAfl3aFHtfAbHSW9SSzkb7HGPiv8uWZzdLKymebRFSgW+4APQn/we
+58Ru1OtSZTdcYE+aaBvjjTbzQsA1L/dEHsH1JDyK9bxtj6hoV8OWHdjnuS3lyAyh6H5vAsF8QNO
SRZ8AxkbQQze4VE2X8xqpzwcItxUpT1ZJfwpYHil6US9gBauydPTyiTTGXhnlTewKyiknLzBcA+4
QzQg4kyZmwUVvMwvt5ZbtTmGN86+R6Fg6ETNYFZgwTmjGiX/pt6/5aD/uEg2IvhF4z0A4PT0fdkw
UYnvgUzMBFEPeLA8fUGgYOZUqMDf6aMeGVVBqNtF2U0920AphWhs7rbtdAdvtNQoWtguzo07ANqB
31J8m0GCSjZmQufqgMTSSsUZaephOe641m2ZN8nNfivkdsGnjrIyLpgMfy/siyoAqkIbZvH4dbrn
I0WwhVmQF0wFrl9ktR0k1tED3pYqjAutlx6zxhwrEHA6wQh6T3WhcIEQhn7TNn1Q4x0b9hgprndw
romWNIA1CJd+KDQ5f05HiCj4DLkGwR6qWimdOSO8SZYjqgxWW9R0VXC9Qy/ZTUNCTp3H8mFy5i3C
D0Dt96iFvLX6Xw2VJTgurMBDAOkzsaM9S4X+HfgahoCxfPynpWXHZxmKO76w2hVxGW1UKlkMiYrW
1rkb+mqeLuP8pxL+fSagsUHWsPuImuFZdCprNfJBjFpUnsv0GU9YUWewQGuuqXLuM1zhF32aeWdn
f54XSr7jYVViSh1GHGRQxEAqAvJ2O3EcuLryCArS1NxkyVROfKlYussnM0xfahvtnwEnamV1OAJu
G6/JYjoHdrSL8fh7lm2/YPKQ4EuQ90geTiLjJHAte9mWg6O3LcQiCrf0b5ltGBpA0odukmKZuviD
3Sj+GcAmTSpMS3AJ7ZM1O9dknTyKmYsi4FVR8PnUk23sDxzOI4x+un5E3gMsPsTpUczW5PnZXhGZ
dxJS3PTM4cJyIsKrjRrvb3J1KV1eVb5407UyT/CJufjD7jag/0PgspH3zV3PTFfqZKny9C/eiLzt
+j5eNa1c5Wcfr4qwtcCgU5MqbNnM+p7VUUvqv78w/lb6J/EigsyuP/P/kYpWotEpFIaf99Amu1Rv
s6OtmBN3TuqlQE5G2UXXQY/wBqcGU/iS8rQBWwbqZJep+i8AoTFsP15nBjO2JQzNAHLsqzGYHC00
8vjB/OiLReHaK7vlsouRG4ZVAxMmIAQqQjs/7UvOD7UX1KM3wicgAEtSXGx21flcEn0VZy9B3Cil
fHjDrw3Zy9hRJUn6DzaIK4fB0dd7DTCFL+qHgKs4r5lLWmtFUThR1kpQJRrhQncmJ3EvGPmNxINK
/aVsEPS8bhj+iXeqX8bTK8slAOHlQwG6Aq9SeJ4xeWdKiRGk90r7WDWHe1vQSTtxzF72R/KqYpFc
oUsz0Q4R/0lk8ZqVpe+F7YUfYUZuaL4EySXqfB0qSh04NVg1Wb4BEWdGFMcR2ROU+D6OS6aG2gFt
F7baZxajBy0uGVssOL/XoPCljEJcyC9E44kWhHX/P0IIG/PTeGAGLKmBalAN5tx8xLBrltvXi4ng
TCl4gBTEVWfjPkV1dRFjVfk86aPMzNM4o7QAm9cI9h5ysi482DBrr0gVVXg64Fjx3HE+mQnSY/tY
QZE6GAJe/uhDTgJZbkUcPaeTwYYiWmDhGZrFNLT87O5AQVwIf2Y7IDik2/MGjzeoKnCobRhkEh4j
BzB3HzW9Ghqc8uxDLanm4O7bJha6FNBFgSJgyoyLXMhG/B71LH1/ucjr1/lJpce2X1QS/J8gUEq3
NHRO/ftDJM3B7TNI20igJvW1Jer1+0rDaTbMnlF8pFpbrIck7ge+a8YU8SCPbTmSzIcMOlyCLzDM
cJs65J10rHS4FrntewxZyQBQlZt0XGhqjJ48CjjGtFbQUPSeChY42Et7PRnNydjAieoPdAhtzWgd
C/n9oeOpyBPno20m+q0rBRGOUz0KIz0AAOj5s7HYkuoi06DehGe7+6X85Vb1/L3tineDFEC9bJZ4
3UTJNDL6idMkS/7qnVHykyAgFiNW34bCu+8TWpWiY8FhEOWVasPZCoIUgeiyFdXgKFHsQPFqVFUq
CDB48VGgLHbXpZ8XuPR/FvY5lDoyL6I1pSCxkDSMk6tqUUZ+TI/CFqJN1PAhyFK7ftPV24Dy3xu0
IS4o22bTFe3ZTLzjs4jIFQ7qX8hxq8uAv9Gk2UAEAmyZ6f9ZXSW6MnKy59rYLBdGwfq7D5nkkkkp
fcVMNaos0pkd0OJPEm0lJCn/UmC4i/MPV3Dakd9p3MbGseee+u52ALr3Sb0GHG27Th3ohGErD1ns
ZzcPi02WhM1VYxg/s2KjATI+/WIur3CYGVc9Dchb+UVnz4CmWRVCIE6Kn9H7DyuT+xKmv5YduKeO
lATmUjSDQ50S4fTryei9au0R2G9bgJVLYS50FHluGUScClnna505x5GVZo+Cs+UQhBJiFF72bNCN
NL5omQfAVJJ/XwndnBhBwXuOqaHC3GxpkIAy05N+qEN4kr2WKizPSJtoaP095/dX+zQCTBdIZKBR
PN+a3BYpUzzoJNYhMHbu6kfU9L4jkV9Ibr+TmJU/Z75iKHgvnrk5OtjhSt5QT0boODoEGkFiZ9br
0vhLtc7kIIK2fKR7tNQxdQIoxo5mMcYLV7Wa0TThiIuLJ1Ar/KzpUrO4XYQehu+vUJQW2rgjTIWg
MH1q/mSxXe9xYzTGlNJSVR6i76LFN8W6WUwjO/x13Fv9qz4l6VQmmkC/7zwluzLisSxouPWxwb14
CrKD9EeKNwZ7gWX3WMImgS74u41YOLEGcNNn371+zPeM6BxySYo3S0HwdX1UMFsXnTGWYbZ4EoXL
lasTNxVHbK50zN7HuLZ4IRekbAFXNEpfoctL4vubNqIq9CS7m/BVJBoeTbfYi7tZrUZfGmGsbyfL
B3KER7IuIW/gb10680XOOk4rVOh6Btxui9sDWj9ckZUZjbviCsfvF7+leizEYBpIsiJ2bsMmA0De
X3WXfsEuFowNC0ZAPb1nvNo5rOUaGr92+HIgn8cRf98f5xW0dwl/mAIPSL2FS8kW+t+rlqB0demS
145Yo2NoeFCTNEmc/uZCIQGWAHNjxDc9I64yUAcjrHBbXU1yw8BAdbvyHblgEMQ9Cc5/1jWvJv+Y
8uxIU5WsSZXWRiAh9otYdqE9ogCShJl/9zvhSKvdectrMujoy3JCs/g9jsiA0F0n3+RRlffZccCe
JD8Jptr184AOYlm94jM3lIQP5pe9oVfJ3I3eks1EE0HI2XOf9+sdqHY+n3IyFjnwo2NYI77Pl+ZN
+ckdi6Dq29pe6a53Z5rmZWsuQo8fm14scVUz3iol61cjYu2iW3GbZiYyV5ZbU+ANViELrEIPV5S+
iW/JQRsLdV8DWyArz547LsGkRwp434+soCE0TyALD+RJTXwycGtpmrUx+C959GmzDy+i0lMS4Xnd
jD4tOr+udvvtTpqp9IC263O8kJnQ0HSp/g/nBlrTH8HvjZxyxzVKA/FjNLI94G5qsuQtZj2g3tde
MstgLBJZTDwwsFPzDby7c8dMggX7YhKeUDDiRPRvEqMyDMW52NJ4EBKyHdUuDIaLRLm7/MIeS1QH
Dw9Ebvwh+HySdg1DlPrRdGZWFn07+E+nGeEgQ+HM5nd8t3Ww+BEkzhyJZUzvzX75b0BkMC05ThdM
4h8XojIeBHr/fZvjn4Y6c3HwAsPnRmWzMxm/JAhvbR3qiSOJyn12kqcBkqNdYfTOJQBZ4r9OBID5
mWffD2x885Xze25JzIfL4JOgRlgj5iUirbg1Infzy7YQxVDBMKb6zAmDzce1l5NMcWl9/7wjXqED
YU/SrZ7K8bHgRls2t04O2O64aTBRkp78TQ8ZOXK/CdmrBkv/ck+E5WCv6KPVrBkONwSVqGPWFNML
Ksnsh+b1cEsEporLf3/GCJ7nn1Qjj4UOQGnXGd4WYaA0zcTqfZ/ZbAyf5fcLOxnDbntyastW4reX
0enejC2wvY8Roc6yoZlgf8OFFrf9OxJuY2GQtkIo9yVxBSzeqT4LUwc1C+JZS9JfjzHIDsH2IP2c
qcHvnN6P3F6TbhMKpbCAqspqiUcpb89nZcuENy6Z/cQaBG5NdWhUVSR8liZvH5YMdqUhjfH3qN3z
6eXs/tcDp8Vbtwug2WnmuCPFBm/efZTF22AK0CWnexFDUjydcO8mCtimmR1IuWlmCEzl0iZovRO2
c1kMFEL/mLuoUnNDxFzjScCsvOgY2X7Dg9NYnmO1sMPqi4FEy/zhumEwmENOxWcmxc/u2CcP123S
1Hq1L/2+mB7ERbQsHzHBJR6Dn1GQT/WTWaNWBBW8OC4825MfgR1I8LkTQ335VQtTmMErImD+OI9K
i7dEVeHtFWYeKX6aTr5yYuFLekiswIF5tJw1YC6hxGl/+TFyn/pQahrLrvf47YNpgn2mH4+w9sud
ckH2FQo8GdL399XtlLN28xQLpMEJec0K10YfZQE7sSJ6QPkvhuo7xGJpF+UIZiNs63b9tFO6RKHS
wmvEYTTQWpcVi702TcjDf9vLqM+61h9Zfy4bT5U9GsRYCO7oxtTJLEOiS3kVFwWYOuv3PlZODMlm
lo6MyAa4EBckD5Z9l8PhmWgZh6mknzDs4tSa55Bns1uoBBW//KsMrUvVrQ+xjhvlpsWZdp6Xb9vX
vW2ttPhgUtAnPJ0vERwCzzWRkdrEUPpIq5ZFgaUVsqER+Ds/baSFSy7rNilgN++ZBeGXcqqMPxeF
3s8wPs7hJaL7aXZnrpl5FbYhRPoZK5NtnMUWdBfkczCHBz+VTCn2xYGoikTLc/gz6qKDiJYCBSTV
m/Tdyl88C785tHAr1HquoXGlcidZCcvnmIrGpssD8hDjfc7FO+t7yIsvx6HRJwGVBmFoJK0ztJ4F
pprubA5tFH/PwiZtHLWpkW5+/KbF2qIX28AhXs5FIZLQSB4tJC3c4Pk8MqbxZ+/Sea55lmod6nlL
lidKxn2Ry6zNSdNmWdpacqJF6VVxWNb44SBOZOqVl25TLnAZxTAwz4mLhaLmnydNx72gT1moCMAG
zL5RfPsN3yQ0nd5/Z7lqCvGTcgX5NYN8flZFR4Ly8t9hKSzgKZTbkIUQqoK5roxGB7TkbBfVgVb7
R/GtXr+bs3ojBO/PvVy+WJjubbzIbZH2jYj2Ld0t4Ic+U1/1KPFTqyOzMs74Wv8HFAtM+iXvkCW9
D7arwFT5AhT9AnZwAPo1/vIzWfRN1qRWcy9uinDy9SON3QdkxcN0so0DDVMFS1F8G7Rq5rz/meEi
DxW6kdyLqpwDL3Z7jI3VU27uabSFLalCpI2A+pV7veoo97kMloyqXhH5PKcicElGhiJlSwCFahPe
Sv+gjHGbFnzJe1LgUYr4p7LIPqzVkguC3nw2+jXpmjSXwhMM6Ipn2wtJv/oeWGCdzzj+urEiiO8g
xYeAg1FpkK6kY8yistQsCLHEgmMzdAXFdxDTHYKYDcfMm/yoIFhekv/vxzgctg4JSHOVqePIRf1A
CYDFYD8BmLsi1iPCOGtbvQT19sG7Vmm9zgXSdA7L6rXuHHwURPCZj9PXv52+2Gje55dMf+QE3G/t
pEYqd6qB89lmQ26qFXPTxcC3xJH3JIiHVK2zlzhflt1yLu2b9ClZVwd7BAvTHRidIjvRX1CMP5PD
N3gYPHmMH1URoNVgaBR/tPq+mJhm4FHOhxIw2ERbyhQ1VgdD1Xkq7TTfdHvUIIPk1euWCk1a6iEr
ZmHRr+AcOOzioHMw/6I/ad/XX4w+qbe5pXRwvfGBdnetBdKcIkg2iAG3dU4bZGH2bTWNJT4+m20t
vIKPFFkDDYLxPqLnjwC8Q+GCKuMLzRmSG/Gooig6JTkiJjmEVafZVsjoeA1xIXw3Q+ovjp1shH1m
MCC4jKeug1HlexIAZVf56FdS3booojAXRj/w6YEqS5WoxhIDmf5wbtVm9QXPx0OEVUhvFOZ473/1
1uC9FhWH4AT2Jz7B9SHWx59tq6h/8uuphaxBz/4ohOrUkcjmtlzEniX1KmwJiQjtp8SV/L10ef5u
DYQZuZidQMY/Q3BujO23ECXg0QZS5iePejaDMNIEHabt635DfUO62yhP4SWoD9HdtpGLWqLKneqp
955t95a5/6y6POL5AkgJp06rQVEH8Vn9165+ERCV5EkWDKG47NNvlZ3MaxYvCid8BDtV2UwgDgZG
KqoMQaINPw8YLMuCZ4NJc7SpwvjQZ4PYYHRL8rok6HGsN+YZL6P1l4wv6xHULJ8ahIQ5YMGmVR94
VGpMs8oqNBC6OJSlROZlRdOQUly3qjsLvlb+F21fYhf/Z+HVbJRKkRVUBqOphBQCqx6P0wx2qEtZ
gZu8+A1PvpEkngIBzzl84CafjhUmuxWWKTxwxkh5mxxK9XBohVRCoal+OwPY099mU0NzkIXSHAUY
/G8V4LP3vAsadOtC1VFQnl2MZVtkAV45EgZoWeCzQ7mEkkRt9NQpdTT8rybTfFIk5Pe2ao3ZLX7g
Fv8aqftb0gpQDfgJhDd2pmzFfr8eFv7pOpSaaJ2jVE9IxpArIUOIHFXR1NH/zd+zX7FvArRF/jRL
ORaSen1Updr4k4fA2O58wbCdC8wTYtnvMLel7G5g/sLx9PAGLvyMVNiYQvjj2seCHVOOmla63JNw
9tRxvcCUT8Axkfi59s0E+zl4bOKa+gF8D0COdOeujgxkCubryRd5gg3pCfb0SjQwaJ7xS3igKt4l
o7BXJw/QovAK2jauT8AaNaHyp4g98+1JgKsoDJG3sneOu8W03crLoqPAmrKKzDJK9zG/im7x958z
2B3JkWcn/H6481EAEBrZVBs9UCOkbV6OjwhLphNVyD2DD1YQszTfXz74Aox0YTGIthafgxX7z2P6
5CF/xXqOd9ffjThNRFvjslgCFoF1hOCnXuBVEg3+s4ygz8ed0vPyr93MLu7srWuEm+whSI2KkCZe
Jr2u5nzkwFPUPM3pJNlwYsVcHQoV3r3RYD9zZdaY29jtLqt22qDDpuze/VD5UeonkpiXA7C5xE52
lWl3yEOiUjxPZwI+t9rFrEJGBFUetTkBE+iHuWwYy/tPFyXvQpMD38yT3NoYstIrPjP3o2rUZUE8
NFDZTZFeFluw+4yKsdTTl39WageorSF4wdos7sKZq9BE/YZuXO++bKRrmuMMQ7VlnjZVV76OS2HJ
na4upiG/l441MEALdCeqFDdK07rmivp9yvb21SJxP0bYpiwUjuUoNypY69mOKGO4L8hPDUw3rUUm
5Z+qh5XodBIDH4U58eE5BQtBYe9DLih+6KLKkbww9lLn93sD6kgPEpYsnrWFy5aJM8Hq68LGlQCI
ZnSBw4id72zR0gS1yL9uI8DGUer/RAXbbNlQlR41fjjaeLD3RcGymtdE4G0PNcXr5ZrBJf2U+slC
xCWcfP3wMhnN0wWI2aVP4TZFSvDJDguZUELFE05E9dHpp8CjeNdryiqEG0zXn1jDlR7hqE4aKtfi
K6E0ZkLlxPBq1oznnb2dtiFweufvCLvDPG/Cq+lcNbM40Gietjjo3CipN8dqGg3CXUIlEQk8n/xu
SgYFiaIyY+aUdrDrxDlAYAV/B9s/GFf5kpSJpKeww85j0v9Q77UWvodPhPGcUGavUe0eSVCUXAKk
fL+DlgIGnXyld5DxTAG6NPMmWD7xYlKV9gzqMR7suCgZWE9DIeFtXUuNbbJNhf9pNwePIv4/bsBq
xyOIGFKyOMSU6ggMlF2gPuDfMAciYvZGyZrvyGKrKneWFw2uL1OKA0McUhul/pVPN0w8yUFliLsa
VaqAZ0/xP9nbA4cpR20ReyKb0KWTnzE1/LOCUF9SPxCAUST3pziA6pvdg6O7FyxkQydGX5BebKMt
LbeEh4swNZa8zXKMNQlqk/1911BR9BsYOBsjAzYaXhQGn0iW9gJIPUepa8ZD5pE1mPkn/LoG083U
02lUmmvFvjT8Qys/WnwCs/OzgJf2RfN5d57eGHVhj8PBn03B0dyJDmC/+2YA9MrtEvyPikuDDe1/
qqBbTmy5WMwLTiF/PM1V3zeCJynMm6B0EwP7sNURGAcUEokdIqr5PbclyahLstuUBnnhOjHr1Ofu
vZ9GT1K+IpEyufsSzajmanO3bPVSdhffrUTeRRDAZESbArZ2xMyOQaPRo7RYPoOIWZpJZ8rPVdSm
73BEf7K2gM974FhE86RXowL7jjRNuBRgFjCGxiHlZg6p9ws6HSGMp+vtOmzKZHU1f4GU+jWbqkh/
EViFIVmZukwn/bWgtoPyR/EKOl1VMYICF8TWGlWuuYYW1okTkN76T6hCR87jY2iSrY4xv6riDO7K
01RZoMNn4jN2qO8fSZO3iJUw29ee2hpfVXtepUTa8MKdbSJaBv1eN7DB9P11fDLD73PE12Pbmktf
8tyjSMfDeOd0jkbJSuNLkyvIPmPgosr8rieDSqg//hjceeVexLokiqvlddTeOOCxKKXvx90p1eym
rcJatI7WhfEE+fOjKgJ5r5X6/CTu77SkW0thM1jbsmXr0lD/O82zeHOJEwC7U48u1NhVySIrrMSj
kto9JhpvIvZvdXLhP4la0iCsNcfRpdQYCuNtBjwjgx+xLgFB71yWI68F0a/F8ch/ljLVTXpC73BN
NV4yJINE9cdYZxbUAkBPwzIWIibN5eCCbVsdEkyURmIlgx78h020/mx9BTstCcoU0CcKWn14scx6
32v2xBHbrdGI5NI+mg5PeJ+j9KZl0u19a61AeheTxSz48HnKrr6PPbkkxCUwswLcLBCAZfQgBYbO
imEKRLrp8x/gP4wTCYLtIFJx2wrWkd/U3ptARAkIrQ+j1SyD7IOU0zHLmzPJy6JVS2kdY4Oa6J6n
cl4+mUxCQ8uLQgsoxkHvpoJ1SDXcQLGqu5/aNvi5idNC9mMMSvczmr6ilBnaQEyRS8ewJbROeSBi
b3Kkh6/vjJP23qrRfTviiXn+7bW1Rzc1TiAnO5Fo595nD23knBsvb2Gbdyc+14WlRmeKW9lAb8eB
HJaysI0cVWUBg0aIli6KTXPCcgyWvT66ntSzrVUjZyF7wl1sZBmn/yppY3taR2w7xo9DAUqq0kWX
IAGwI16tV/egUta+SJgVhN60c8OOLSTpqZaKamWPdiuDW1/5DSvLgNNkfVPpUs6HvVC535JMwHoI
5/5rahnWDmm4S/gjm8jXbdHJDKnBmCK/qcNzBzUAKQAkz++H5ZUFysr/jd4E3P4Gg3X9HXR0pm+T
sE3/HsB+h2sW6cTk9t9Yr5GQ88kU2Dgp0hTmS5OixwPWbAI5UwSuCwG5fLJPDuGdHn+Yqs1+kjCB
9EyPaz2yzznAqfXx003M+2cu0EZhza6O+v0jZC0cAG9iFzTmrMajztn6FcsCOGvNq/j7qBepGNIT
ZgS9PtEM8mSbF2KgNlX+CH5cgHGsp6iFq4P4vSgOGjI7OAPrl2oSJxkbwmgZJBVcBBYeMhPmR/pv
c3pEh3rpz973apQFvvh2EVxHg1Fpy7EVFYinHC4f+N9PH1yG1ce0BZi5pXzA3SWKoSDS8+1oky6T
LmKO6aTXb+ZcAj3eDkxGX6yGRtdwUfjT9gxuwCdOnaF1ViETk5j6gDwfrh7YQsNeG0pkGFvw2+EA
reIs+/mSbm/YdHYxQeJhNTDIaxDKHuuOQG8hqE431lPIzz1QWipg6RslMeP2N33qWmmIxDV/n5V0
H4uYwbpIV+Digqq/UCobAhR2Tj+nv85wjllxBnR7L5TO4PlUtg7kP8oWW2GkMK4TVae6xkUricWF
tBCk+d3WZqWTKB5J6t2L/DjVdJWyNYXsQavwF7P3teN5RQ/DZqIWf8Rm1McBXDDK8NjxSLKcltU9
k1pB4Fa/Go/VY3B/04ip0Anzofqtqyh+Y58uqt82qDuVcc70X5whyDXP8rfHDIPbAKzfeH2ctdrd
ObAOJOu5XUJeDEs78zUl6SgaptmbF3YCe2NeYs4bu47KxPasIH6ew/TAw3kWLN8sXQM/GhSKSTBY
KsPrfbedSeO0I6Yjuyu3+ryeAfzZvO/DaCkexrJUpdrAmJmKXe+7+eJVs2k4mz6c3N36w9SWCjwk
6UGx5rfnLpo3gZlSSIoGGCmHZEmrj3SnZYw7cFYVVERQNXgazbQvCrItPvd3VMInuActPKoB0yeb
oGk/RuMaeluE/0j+YQdS/7MQy+o/EHInfBedoClztufT7SEs0WYXBkVcQnIAuAMZzm9PIw+eMLxR
SR2LgQlsmVm5RwhJf076Jw/hLO7i0DuvI3EKoVgvfmd2+AttS5tAUJ07GDW5zeiZWxg1ZjuJ7pbN
2inRrm20mOiu4fNb6ZN32kjldCviQvmZ/FZPLZrLo4e8/SjTk6jHJzdP8BId8cFrn+Me6aCR6xhx
h6RmtJIMXuEcuXBdUt/H7qPVWbWheVMsy5ANW3gx2mlCWFGoOIH03hV2eYF26CZDDvkK3UK4Etn9
PpToMraBWg+cOWS1HXYflOhrzSObQYV2gTC2fS+J/NeK91sAQTDq4i9nTFeAylxKWsvpSCdHtKO6
Opiaj5WziHkn8KiMALCfJyqdtNUtZ4m20/uTccIIhdzNrP1rokIPVkFPtY5c2tw33TjMc/B/FqZy
iXkXmpzx9VIjlueXYS+chZOe7gpjD/qCsBEE7hFSYA1bMWEBeMS50SjAoa6nc5AXzBJj5B9sV29h
28TgKGj8BfSvVpfb8qRPefxetJjR2gUe6VNJtOpt/+f8+b5JfLo8MOgysAhOpSN9bTg9WQqpY5fO
ntanqqj8YXDa38W2uZWlrdblSESnrpsYZZ0buJ2MPhXMC98vCWKa/+P8KYamlCyVpFddj6lIivon
pSOF+kX/5l6m3kYt1rQHE3lAUg3nj0NBKjb2oSRKHuG0tvMJ2vFi85/JFJI3ZZmRsmAjYCWDg8TQ
ZGnXuJ7MaQf1VBKqPVtd6nzwozC2Ki+WHcM4ZHsD6skMHStBSJ7gTmHgZmBp75VYX1V6a2TIXEMZ
qhRy7qDXalCdWetMYAlEcjX+HW+iwPrro6Wua8CMBQIdnPLvzcyEJ8imMKFL0AvcgcvIs2UdMXiG
2/9prjeJ6Sl6fG/0nUDHY288mTFfnFnZNc2UFtdWPr7GA7i8mJ30SkL746m5UOH5MYjRqo31QSet
Goo37N/0Ap5DcrJYxVU8P1lo7Wqn5gRj4gYAZmUIXXgYUXhuO1FyYGJs37TldlGLpzqwWgXNUC8d
ZmI1NT4Yu1lXXG3eGLoKy9HPBlatZB9mVn6xGuXdcO5KRj9Y8hPShvkYT2ZyKdDueZam30L7KzD/
igwEcWI0Mp8Kuh6YxItau+9rV8KlS4ncmqul2A5Yun2ofkx6rw5DZ9rc4Hmmus9gcRc6INYXwGkZ
I6nJZC7YZr7Upb9SqBDMNl+/VXSaiyijZtoeNCA49QrIvigMPrxoO7s1t2XSSPAyZWp5RL8rBMcB
JYkpTUolTbND9p1RbFLYcju8q7/mfwmf3vsTIxDwJMgizHz0KlcraxnSFvqqYRMGCpmAIjgBpFkc
4j3RsbbBHepqGtNpz/wnxQ2W7GbiLz7jTFedLjrVVDEtEyCmJmv9rMtghRNoxjCDtHA0OhSym+Sr
gfR5O97/iVxaVg1+C4XhtkUMVT7Xn13XuJ4Av2GM7yuWA/nnOMxFou5VzOx7u7evbQ9Co98xphPs
mrQbiwWm+MZRWSUefeuCAH69x30oL4iOp4NlnAVFt6Cdj8PsTKY6c/r33hPPAxZWOwBToBhfxCXy
l7v6QY/EIzCEr+eAttIw6BxOPbbLsAUjOvDXjeEURpR7yX7me0WaXSwo0eVqma7jL9c/O1GqAJln
cnhLTUdVUyLe63NN/VsMbHG/DCur899YD08t5CJhDRuNrb8IMQaNDBiG7+QSf0M8PWi0RXk4fVn9
fgYj/MvRY/UkOJrTcbiscZiXceEfHGQ4wnA2ksi4g10n/7dhLRPdLJyccL1z1lzJ2cQ8KrYHvsDY
pPSzOrH66Gzv2LZOpX2SFqnQfxDXwIReoeV3rXK7wu77QhA8EDRRzCNDb7X0uycJrDrnp15+AChn
XbzQHN5qGSy29FKAN6Z9zU0V2iJSiEepqmtGJWrBR5QNB3TV1ABJF5Su3pkwFPLnv5vRwWSFp9cA
9lrl9m5iT0pqKzM2YdSZ1luqbLAXz/o/WUU/DI8zuXAcjYr9Kp7WeLsiHtW3FGH0htRRVtzAakT7
DwuztQKZnf62yBV16qi+6Eb4d2UyfhmtS/4RUifPnBumwcziCEnO/2ZDaRWLOY7uFt6kv/7Ue/jt
YgNoWeMoRCjAeuReMnbqZox/L0+VVr64F1t8+K7sZfPKH4pLiVfmfdbj7raQ1iyQQsOY6+fHeTRn
lrEc2LYcQhFPU3WqryNfHxAfyYfII6QIGdeVH4g+wgEpYi/PdFzqjrj+hFAx7wPlQ6YFYb9Kub04
nT+gjQX7RxNpm8rpzJuWedgIwT19E08ARZVVCFsYPx/lSCOVsyFd4tgFxYYgtX5h+POh3RsSlAIJ
9PvLWe1Q+XuVEH8nl668YuqLwPT7N+SiJlEIEtD3Vb9FDFImmCTOVHEKu0GiNwr90K/BQ4AmxGNr
Soh5SZhc+qxrqMHxTYCRcWPDlLnDu9oz1WdE1cEjThJkoFUuh4Nn5Xkep2kKU6jS3fjrm1eoy6xx
WOC38LgpWJCMYdBWMd8lfjuz6HknS4oMDObA/cfBJYiJVGk01jwCbvFd12mut3RzU1IcqD4fyPsK
svEoseYJdcjSQebbowR3EC1z3RqtmBNN98d+9ycBWoxBF9kP1pvFC0Z3i0n+KMU2fIoomPPbLyk9
AQpXuGaMg/jNa6seOxk0GkNINie2YPkRucMbf/Q6mnWydM9IIHkRg8vDx8RoYjIDD+wZuvm7EE8R
7+tphBIdgWuNwPk1QAb5GmASgkKvzaUKv0EHXfGcFkpN+Y5KcqjDPcIfSHNqki9E2kyoRXk1kGtB
BLU2djeBSmdWSfJOCrZBnZcMkbLVX1UExj9mDSFrWbaq3ENR3fi0NkTZBm7qvN5g2Wy2/9cJd/LR
t9r/CNGa/KXF9DD6xox3opOpTsIJ3V6a4bLEN8PjPO1uzsthD/gPDLJn6LMSPDHErRiPQebsQjXI
VSrjh1O7QXs7bcXYHO6N+/O7ZwX9gQnBkPwhtOG5LhaD172BcFZYtcXfM+UUS40tUAmBWGLaWYij
0+Un9IKqhgW5+WTu/ufu9IcBRuKVj409xK9k9It2OPvcdmHc8ThStsOCMZDKl/Hc4bVvvVAliF9t
9YAdAUdg3mdRAPWhhxZp/sbXWuBpB4yGt4kUjeM6eHH5U5PT8iqlOybAfd6YfWHxz4/KejnSq0mn
9vVNsKSxDK+KqetXk1FKAfFPcFjczb+aD94h6jTz9XEBs444pP7C0EL8EcazBzZWaDU4qRv4s06/
B7HdikQfa+S8VE9JW3Nebq7m5UjgHYwpVm+xUJZJwqKXJXe/9V59xhUZcPalKpWdpS5hYjqku9eh
WCpUZoiwWYalUcxA1IUnMwhYjvCbfGuTGjvVq/zXiIbKwZHqaGIafPJMhjYHoR6UFv/oaXQHBuP9
K/NFoAhT6n5vgdCamgvG17f7FMfNJh1QMpZwTaiO2CM5trkUKTzcq0I6B41EEX9ya+OuVc8Y4CE0
5gbjfBaQAGqAQ8STEGi2uGzq4NBRRALGRs/oXGJ9RDnoGWcXf4yFndR+D9sJV/jUA5h6NNLLDL1R
c7/8uH6XxdG38s9vJ1a6n1aqTebBsCXidP6aB1uhplpmUqGIxNdnqAlH9R+oGN/nrqlXjuVzbiNJ
7iMqPAa8r998qM4pJWkSjPwr2m6LGwaVOpseMIIpi6edg2P/fT3TKglCwE2zejtptQCEYLsmdZCC
k3a1RYkCIw97wX8A1F9iuWdxOpSiSGdbnbt9FPTMFBURoo1w4PUZqHH8nXDNa6ZDV9K6S44keyxI
imjzu+FoibiK6b0P+Ks4QvlwkNg5coGXzzEcbXQic/D2PK4RVVvYa6j/ANbo3yVFBBz4iPmr5W6z
og+ViCKmDwDyIu1kxZTgE4X0j9Ozje6Bea2wV3k7fSQGVk9FhFTbBfo4C+xPDPN7vA10yG1TCnDB
EQJ6Qq4Iw4pCm85a1zeE/wD8GCHYYZTekSGLbNMPe/HwFdNCPyizn0ABWbUS4YmOJiyRUMdjL9oK
/WA4XbXdu9vvDbbCeLPZOXZwj06j4n/Isp25LuiLi6YgFujJGfjqaZ8fZj9kiPQumQbZaAh+05nS
MmGTdD8fXcO1n8KWpyComufjiXMG+nMxH4u/wad8GHGp2lCeGIu5ue+YGub2pipHtqLOf8nIFAue
eols9QKMZBlBnYhrdv9AMNUGRoNQHLgkWlr5VK0JeHn7mPgVT4bVvXrYZ6lD2Gg4+G1t8Fe9hUlG
CPJ1Z5y1x2aQbuo1bte0uhnO27C1D1O6MBlnvjhzm8x6Hg0lTXzIJuM94XHCR0WhvsRiyDpKXAvl
HI0pN7DrncwT8mYQdhvi/AIA4l6lhu38EeUZ1OUNSQpX+5nrki67oQf71ijodXAKeooJL78Ivhbf
86Qhl98pi78SR8zijBFKHQsm8/SfQsSKcBwggWr95gbzAwOKAAahVn3h5v+ICVml15rODZc6Ngg5
LUrSZ1wJacTVCfqVib6ksVJRq6LNpw6qce9wNG3G8R+hCLIYJp0zuGX+VQjdfqC+bdYXO01WxShm
/KgIgOZ+sC8yif231Kcv9jJLAtDdaZ/W7nJdzqHAGXglfsj0VECjq1SNAz5xxZwsQfdFz8WUPcYn
2x+vXDHrlZMx3XX6UIyxLmW1qbUPUDJ2zwaBqgeDadY+FhucA+4EcnMRMlGfdl9Xf19f0C+gl/+b
HSvKcun3IfAUGS9ZjRQexdTJ8ZVBUHlteuPiZ/yi0+rk0SrrKykvms5idcnvU6dm2xTU9dKIqQ4Y
MD/G9VNElEWVBP8DaA258Anhn0zENz3cpt0mLiN4eALx4DM1fL6Job5tex67uJGcbuzbq1ZaOK4U
EWftS8DerXglrpLKaxjsrgGEOBlv9WiLPlLOoLWjEf0Dq7CUbCVxoZwe0XDXOdemBdwT2ZV/1juA
f4AH5/i2u2/bKFI9vtruPNGYKeYurZBiagdh4TSBYvBNhhrSVR1cLPXNPbW9aj64h/Y66mOdFqYQ
g3OH6ESOahnC8xHnpAWL0WvLsh+S3h3QmTv04JB2PxqpQo7w9A8iVj9iRDdoToT8Qm2No1BdW8Q1
quUfKIkO/u1NU6FF5iKkfjeCytrgNxHWgB9xVw32va0DR39iFeO8adKDsBSNSQO6JTTBsf3y/Q8d
y5J5ebnzSvbt3AynyBrRiwsn9wdab0/TEJGFUvbiJ4WIayBUwMvED2X+QqG6Q2mfwEA6C05jXFsE
EuAr5l7+65+du7nqjTEgArwThgGFJu1X0torm0+3nmHQ/5kCKQy6pX7cKkbChavmarppx7kZxxeQ
cKBhLmB6HBAqNzAbDsRrinxgj5aPzVrvU45TQ6E4qsKZ+dyRAoLguz8NWDtQtnJ1rZCE8P1lNY4s
eZD/TlRahz4xvWWXIlywB8UWWWv8sJP/tmvhtxgH7glhvz4ZdxurOiFvChq+LoSAvNQnVpO+pHJR
wXnp+q9JAM1c0bABs+1LdPYq48TdlibY8YvBjs/lNJ+VyKHO1s10xt3anmGnZl9MpN6Ea23LTvba
8wJCewHUQZhPXJN72QD+pj0lBnyn41NGcCopMcMhynmUcxlsgzbHVB5lqW88xItlgaqbUxBpbQo8
R15J7BT5k/jO6B24bMSS1GzIbO6u3StYgl87z9AMRXUL/QibROITkrUMcF0BPNlpM0bevnmLZCWY
yva4lMCn7aKIUdLuXNSZIN5LbBKWVcl0RpLtagvcbeUhUqE6KlNgmr/5X6vX9FixZrAqwa16oH8Z
VfX3E9ro397m3SD6kM/yR5rcThcIMDkuA1XALlKKLzJKcW+JTL7QEbfTbSKAjd5i+VhqFIFzZflu
QfZOBKyxUrlAtJBPaHp0uEfBaTnLh8ceyiI9FRvx0K+tRE7xbUHFd+Q6RGT5XEm/uempw4Cy8b3M
vmV9sXjqHNdXGP0Vj2bHneMm0kRn7Zg+RwqYD3BV14SYmN3Jl9UCe31+KIBcrOeGLrc09aqNc6+S
QtSZuAWzSSocJqv+izMV7PO5yljuX8Fdb63u1yvYp+Yjgjb611ZEmMdoKsTGf3TeFiWzrmGyVLWk
nrHInL7b1lFEFcsgmhe8FS8PqFLdyuofaiLezVloAB9nrxhq9JtPKTQBTzI6tI6dDjg3ZZPFxavq
zSWcPrii6lqdYt4dOfFE8gmxdyQVH/UV4jOAQOflcpISYUtREm1RcC7SfgMll+o2HNAvtfL4ig6k
BMN+UHcVtbB2TgCbrsR0blIT/iKNOM9wQgj3booTEdOGqWfpvoAYN2KaEbfNHWf3qXC4iEmVXEiE
WdHnmMXvpmzIkRfWwIe0Qog1Q898fYli84Tdum0vhqAESP/lpinwiPINkfbAKtLE4ySQnxQU1nYF
VzcGp5oUTPaHq/bhoLEcc2XqPItAPv06S7tsyU5X9Vqm9X5f6mMoL1zbCBs0z6FwrqFKMERdBfol
8rUuDuGOLMx7zANGUXlx7hQkogidZB6XK4pnYMvWgfgrujcYxJhQf7PdZsYgbPOuvYQqpVUrqAmQ
nE5FRTLt61VLMAhGGMqk3vjsEE46/YWgb6cRrhH3PuEVwkwKq071IFLGcjFav6KYywbuqtJfJe9C
mD/tg7r2XB96+cT4fdN6ttkX9xmxb15RLrbxIOhmCrOrGM6Yf3522Gn/H43MANcyRb9AnVwe1+ku
WVLy3CRhbsx2E5oUhd4IHZXFBJfImIBZ308QkPVxI2DXBAf5ipUNPbn96URldzYupOKfxmsPhe4Y
gaIx0XSpol4GQHfWHiVx5qN38BB4kqVhKYB56FsH+mOKxfQ6nP+xr7Ais0wE6kGggxUNI4o63eiW
/GfYgvhMdxq64x61eoz7V66zrkyBGKexU5g8qoSQcxzFlBn6XgI4u4bJkEOCEeWASK/GkwZZKrN6
IPZZEcxu9YvqoMRRoI3T8v73Mahqa6ZkE8hzhPlwmiUvT3c7h+NXf9b/sYdQqSJ+SKLy4gMuOhTJ
QpRwVBwUS5Hf0PLpYuKwnMsH8opFCbZxWkYAtkQo5uOn4xgfPEvngeWmEIGegNEWEo1ONvX7Q9vE
/2Ms1Mn/VeqD5RHGSoKkDuoQuoQQIc209l3GtqMuExDoEQ3ecJt6F4eadhT2leneOJ/7lr/gB4jz
pNV+pfskEK31AcfAfgHKFnHt1xF7XtPMajSztOle9cd1owRI3X2GHv26Px7Js1pTEKKoThasRne7
2KKO+xzg7lMMciQ6pyn0rmAyEP9qbEBsUKNVFgwCwB95hdrIrIPT0M3e46uZJH3rveXv1UieXi/R
rbmtiYlximFbpY2+KEV7whguTOojM005Ph/SGk1cT/bvOizC64dcVkftSlbNyrBTuBSx9pLjKCB8
h7QFwMIW+hdjrQgtpdTmwdKDAS4WiAlfY5pHe61CW+VYmCtiyYvRToVDEeXGOPWW23F2Evw6zhpf
sY8CNMpo3NiV1DqHwt331fRrfouWdOrftKFixthxf8SW+d14NSYGZTNWO6D5PdtB/AOpoaXkz8Xp
UuoX8jt3hQvMAEDnnEI8+MgUctCggMj1ZYhaN/YDgksWghfpwZLo5Cx6csFp4j2iRrt9+j8Q7sF9
H2HeF4St49kXzxRt2nyyggxW9h3qmYwQbC3KSHueZ9d2ltD7UYCXrv/RSrcrtGx2acNVytL8UJ6x
y40Mn/LGycc5qjqDAxFdF2J8doaCoNMTsbDZnwKDyH0ArukLBymAFwobTXhpxkNjDq4Tlr+aa1FP
isbeeIDJ3UD2OKTH7KNvzsVRnLTIPMzKUoTzVtY6BRGOp3wpr3ej+iv7nBvRr/pfnA5xLmcEfjPn
jwJqD9PQdH44gnCMb3JTp3zpyAYwL9qY3Zbn8A8H9UOFBpVELKxcXX3Ob7I6X+f4GHgz6GbGQ3x6
j38RAeekKNA7/CwTMbAblL8mk1hprSSVcdMfKwxFd2qdWl/TUQ5eORfQwEkzk+lnSsae1miTmOBu
DgkebUtFvgkj5yBXS4FGq/jm3x3Si6fkar5X2Y2zIjXTUGfVkpb1B6Hcn1Oq7V5WSQJBanrF5qOF
jatkr/SmzFH7ob4SlVJ3s4ij4mKHwNnWdXki5UDttvju117klXUlrrBA3ivw8e7f/mk9+wYQ2tkm
VtxNSWLQoccGxDDvjJaMdGGibijfBRi5YmrbP/hA+51FS1WWUp6Y3IsXL8h6jdo1TUaruPGuPYXI
jlQRgiNLqss3UA/mLZiS0684EovvocITucGpTrhTDcRnozfVGMTZw4rYdaKw0eVlmvHjRBm3Qo6g
AuGowTls5HPezWKM4ofRQdzBtuVrgLJvTDQlWF4X4LFAy13a0lRP3KsmLWRS6yQM6VaFSSBuMilL
XE5uohVio2B2VO/UQ06/2B9sJnggknZwDHjJUHwA+f30ANd8JmSaOslUFrD269ggyeMPpEH9Y40v
ljaqyat6n8OJEXQ8ebtaWtVyj0OOuuag3/10NFJOOmhfvtmtqhkAvGmlR6yEaAht8YQMaIE+638m
DvTz1KWRVTvrGclZBS7qPXeMP96pqOL2dB9RIDr7TqNnDql3hJs67gvg459DUDd2gPoUY8onVkaO
seTj7+no5D4RIuI2Og+Ax6LNxTFb1PMB5culfSnGBzlq6bwzAE9ZWPaPMeE2KCZQRkCutT3QYZyf
czabiy+JLE8BF2VkbQ42xApLCBEIL4LLcZ6UmL8J2mqT88X08c9g2ARNqZF29Qs/0N3Hui/v6E1Y
IqQtQeOzFfGBae4gdB1b7qP0kdW6h/sWQQx4yeoXXbz6/wNLld+varzHFBWave6UxP9IwjuHS+34
YyHd01PSKTonKG9zjLM30tVPqqOU/iAJizXm5B6QP8VR03fEUwjeBmQSKVbAVtA1m4dG+cFYjk5o
CSY0sL9gaFWgFRLPpHBgPplfuYasKLHYyodwAczlDtmbHmkY55xbIYAa0wsTc2TGYUtczU0eU+RD
fCr6m0PZZyb8V5R/FFZGObNdAgZSFuBOsk1f5G3sRt1CjhpcQobVw+1S7EtWOyqN4Cq4+dybQdSH
tkMpHR0695WGt8G95B39MlYqOfq0OiAl4PIsX6+R9WXHJYBxo9lCbPRcULzhOy5NZGfZIdsrWe9e
NUEvrkoULqL7NXzapCu7dvcYto05YW0H+04CT0HMrOi+C2fAwMR+5YehdyduaLPi8EWK8YmiyvSa
LMLBFyiAHXEtJl0NO8Z66dCEOfBrRgKRtHfXMqRoG933ZLour/w2R7clH5Uc9TYO6n5Z4/HGpw1P
JaProZOJXKRPwaraYAHyWukxvAgT/mDfevwoO29aPSZeZPHSOeFdvbbU5Vwu56POA2msCLNeFbhC
DH4xaW6czJ+mvj7/lmB2tyXTLVuXjIaItNvti/4dqA/NfNeydamQFb8+Xr6AurgMKFMADwhWS4Gq
/d7aJ+zOq0Wec3zRuG2C1veFI4bXb/lIhFvjiqk55fOQo3BhDzGjwAL8pg++wXpZ6ObIpyF2R06G
HMQITKZbdcNbTi2IKC02IwSh15+0Z0/5rO952s1g0seOMLjV6x6XZEhrEPn5vFZwjLEUVYCrLnKX
f6NC1US7O3NV5XukRmphfNkj9tI+b3r8USKE7DbRi3xDRTpOmPbSSvYSkdAiAh+X7T7fW6SlgY7r
oe3TU1jC5gj7+15aidKlscrYwOWNg1YyaAX+wcZPTcsvgsNdI3l7tSarzhIuRCNwCM9f46H8+Rd+
tkX5HV5OJC3m7WiFp06AlOYUHEjgMvrmNdO6uQOCHzZcvb1QS2I+ADkGXtn7HYR3tDjMB3WH/djm
HwXIti2wU3Po9wE7c7xVbTJPuhhbfZwvgzWtzA7vthypKX1yMMLGQss3f22hs1uPrjN1Pfgw2HJi
5jS+3My8cvGmxmJ+rFheVaKTaK3hgVUuvl3UQVvaoM1UmgVvTj2pb5elR3CFec74zWo36Z6Krega
iiIwqDawW7jQVxWDw0p0PaTpWAdR+mOetX05DqAcJ1+++WVjOxGHvAUUIIRW75cDxqKXpVTx8gJc
xkFhVHEGH0bBSphdQIBK4plhWG6SZ9hJw+Cw7yvn54yY0A4VzLUEOd/yL86/DdJtbBO7dXxIzyrF
bUBDC9FtslBNwgQSIRJrqsgnnzbFEWbcyuDUUqaz+IVywcBS7RQOJItLsvzSQaLpE11yxMmH+RGd
SR/GpqkSxlBPc/1qs67T6VxGrtUPRscPmsNtEyToed3rECQPTg/m974dpc8ll5VRSqv1EaivnWVz
SCNR/sxn3C+T8VmrH0M9n8e09tLVQpkdh/7zfl98LvuNSDZaQ6t2yiQvNccq+rYci2CTHu+DiaG7
M7FQw485k/QJilyLlG3fCwZ0YuxeGfrQLiDSXzz9HWJCVPr27Q0aV85LgeVj6dhEf1sRX5SjGJH5
wMToTqHcIGybDmPOA0DKZpaKsu/xHZ9z6JxFegzHfOBxwN4tF2y60At0CrD7tu7BNWgDZSPauik0
C6p9G1E8VSrbe9dWku2aJcVvyOdyXgvXmAMQN8EGD/uGo1NwFKjMhlIoI3fA6rhtuc/vKOfCUsDm
dfkHkO5WI9KR/8GD98ywL71M2qcbf9mUaVupFAJNC2swTviFAdEcA+SdIwGd1PgPZERLR9U/tgaW
7d7tnswsZwuUgVcReitxH6uH50BI49QUDfhEaJprKOwepFFg7XMlnJb/h2r/U9metr93YmzTeLzA
xLggcx7lxVcoHcpvn6dCt2ss8RXsnRxuCoY5yP4dSgsOEAh0Uwes5YQIJWXwxWgyG/NHW8JRYbT+
ZQWYoQrGzWv64e6Y4WdBKVSvWyVMvI4GKsHOSa2u1bZxWpz7d0a8mYtiImHszGpkRVxtbADwpe8a
uEtOsq3ufU9zVQHU0hb6uQv43qacOXc7h0HYQ8Hls+1hCGkwERuBWjUY9UYbBqTqbkjvVSXBfj7y
GCJD2KuvZGTnPHTF8l9yKkEghkmZdoXuMA1c+Ro7rXbaBppOqpHV81HGHdwSpWZ3jFNCb/ruZz3I
dABj6pIglGtGDKdnOVknEb1wkLrlJ3WGztBAIWLLiaVl5/QtDmsIRKqgRL5Zu7tWTUB1Rc4jQ/zN
XmeAdJD/vuTZRxPEPns9lKeHvq6Ldubh5/2mrzWuesNGLigJ9Xhwb1l1/gvtHmDz0ZqdrsT5azel
QnCy1UkItWqMimewB8dvF6LvhgBQKtxB7i1ua84XFaKpYuAD40stHiGGC9+mEh3HX3F73ehfQVmj
JpMHIjsiauRSZBQ82OybLLH9D3EXlyeOQwlvf5OCrYVRdSoBkdmgeoAGmAxfLTCOOyDkvuw/pzen
0OcbTa50XRIPfcnJXU/uxLK+bt1uiN/AyRdMWAb4Yso5ICt8NRjuPJU+fPzTPCwIGeGn2r0xrhs9
hOKuwJrRpdX9u8wAgrIU0s/QkkJ+0gw7cmLrDw2Va4bnSgPAYXkT0yRpwhiMNmD0R28T5GyEU39T
Omc+NlDmKSxJMKoxsBusgIM950hTkPCQZ20k4+Im77PzVI+tuRHiF8jtfiJ/gNDcibz9NrLkKknb
SeYHn2Yl5CeWIygAOAO1ZuUkKHNWIrW42BeeDtzDlRhTZlc13ED3Bv6UwwIGQsz5od0vVmwh37bI
fMIUn/fzwgrYDreB/Pi8ObceAM9OdRC5eQvvyu1YUC2fXbtPnWGbLjuUl0mZmWaH7ZC1n36wLx0h
jfFOrVUvaz/sp3KiOP2fBo26cj/EvRgTw5xTSC2Iiv6YTjmS3L4GgCVMv1UWDMqL4Hrqi45A0sqZ
O1kmuPUm7LAeZzoNL5HGVD+PYEZnHkQyxRJCv7aTWrdRzZlj6q7VFAgY7AnCQtNlDitJxlQkawEi
nBDTMWdOqFJBTahQB//W6nUt6iBF2mg5grGOcNmQvo7FXHyXYICV/aTWhWEaEJCPsJuIjrA2NKph
ojnG0O/tJLi5fAjHUqZjvCmY0GZA+DqZ7OyO/MYfONcKhJcrCsAl6hSoX8FLwbfsBlEB/dfixBNu
4bZhBHcLNlMXDUsHg31v27zU5VWV7FrF/p32mATguZHjhuKQTXomStpCXsFDntHJavH1/gzMiKWf
PLRF5KngNji4RMpTIdXskblU4Y+4jkf9uKP24V3R4UhERCB2YAPZkfkMlFtyNqwdFTViqLA8ufpQ
ddEIV8MuqYL/fFULAGO0FYRASbdL5Q3p0bKrR8Wkeu/ypSq46yijKa8R2u4KIDIfWuvOBpnzoEFw
IiP+cOANZsIvzrRcsYbJpePN2bGbDfgpoKqvEFQxhLwY9pWC/S3EgrpB5R2hhGKVILzxd7Hc3gD3
h1vvBV4HOBptUr8/yceLx8Lcnx/qj31gEgTX2/jD/C69iKT4l4uoc4BX2/B2Q/hBTPRjfhKbzKsr
kvGLCaRCSgl7xwD2PZhjZ5NsxYEl75CntAZtC/o6nRP8TXlbrFcn6U41t/nXof6q29ZoVOdI/Jvp
Pd1sa1xnE/BR78NrNPSWbrnOkZi/ZIb8mqss/yQMkiHDI0CrypaECjj309f5KwDXrLiafj+ZI08O
KIdmjDHTqw4naqZJ0q7RBSNXPfS2ZURODj18BOeHMxXr7IZorrGtrJDOyKi2u0M6/5I0JEYJHKS6
GMLxvaTnLfP/ENFR2ML6tiNQRBT4zWLe8r6+HC5G5Yi8nZUX9ilwgiQR3odZLgrY0BGtR8OooXNP
fr00piWvtwV8eC3uCSAgaMz/nKRW3nNMdAbjbHDvZyVdmHMBo/++CAYHbLnWGt07e0r10PGFy0LL
M9abezsPiGKCsW+r38SNqLdpbIZGZ8XXOK2CRXcSv2BjY/GyxDK/nJ7ab7wGYQrJNq0ffoV9jtRJ
B6mmsD25t0PZiA/hD6GTFFpIKJD/EHBkq5ZR01wohzfWQM16T9pwKSO/XY+bluGBnYprgoVKeYpo
emCrI9sM5TsSTr1LUv/exUrqEgNPNFuQ89bQBX1XxRVgMco4C99daz85ruSvGKBPiIUavx9vtDi3
du2xP5jcq8ZIxWwtkngsFm9CVPoHWuo9NecMvqA5YHeKVdVnB+UbrQUZdkiPTaegTB2hImu3Z205
tT+Eckf1QuAMXZpA98ivfWFZM6qDm3APpGcpP+rvWcSuytL6GAPtF7H4JGFvd+93qXyWHigemLc7
agHreLRFZCPuFm1EoqOfpyesrwSGfgsD/i85RhXFRtO1b8VpYlVHXs/tYlHViTsPFennupx+SkL6
f9dWije8f7Sx1OJTLXXK1RfIjKMLXqvwubKENKJA5WJrd3uvyGapMFtVs5oTtBURpKzfqS7CZRs2
WBtzxpS2mlFwDtJraHVBCFB0JsltDlKfUuF9xgAudDzjZ/oy7T4t+rFhSAxCjabFBjHPCGDYt5JL
BoWuUAKkPxaEZhuPq7Hot3kqywtdaCQSoAh4hUu4725j6crcKHCqeQh86YBz/6FpRj+eSesmBz0H
vZUTIYfOLTwIUCaphdyWHYoMe2ithcFy/qF/kUq3EFLXcXSsRwLFd5LLkmkpZAZBSbwbLh0KoEkS
PLxFEDNVaajozgEUCzIVoUGaPs6uf/dePl0wrxLVSvHT9hHRmKu2EfqtBDNwUichFmHe60IJOopx
Fomqqr5K2abFZiYrG/aB8LutCmxgx0e5V3lQGf8fTCgtzQGKK910qdj4FyqvgyA4k4pMm0O6O2ZW
HTtyBAotlZ8n/JId2Nlna/ecw9ZjMSAZLyBVBv7Ap5HorqTSJW1d7SFknXcF7Ira46r6S+tOvEOE
g5nBXtHYc7CSJyInaHGPruZtRPabIQTUsanz401WYdZjsBHru8t404F4rZ624BbxQZpTO49RbQi4
qfy4WlYTwrLPC4v7yjnSG6zLmqarZmU30sdczRNYSvbdhWgGT0sLbllJLZR9QLzkI7t/S85l99aB
eDWifXDSnUl3eJOBJXO8pfuDZN3sFlWc5dL7KylvWV8pPO36eQojgJeRHeFpGiABDEKH3XoLkeNB
jfDX8HvRGM7v5juEtQWR8FA8K6NByzbmWkT32gi63mq7aDdA9fKeEI7LAk3+Z0O1dpdaQ2qcD/ry
+IFwSPS27layjaopMaMfP3xs/nVWGxs63qsD0qFoBHjq0PRhmzjqThLwRcb1eIaOrGPElAmEY7de
ymZetjw2HTrHQ6wt5KSLtRTAyjShibmAX3EKwxISHNW8+m3hREZgSd93m2UB9btZsY7pzmEeSimZ
Jifa9RauX6hGHQYz6TC5M1nwckLk2LX9oNNXhydPIr9RqCglcYqIx2EpJJs6UsbkquNYjHFmcmju
3ruuSvmy/il2K7uc+5cnIBHrhv/whQErWtq+ZoxJj3MFa+qKRP0iu/r2r8FnXLhtjZhyx04OvheE
mdOQNXlfzNYRpvVSgFEvvszgVaQ+9scSrX7g3IhUCglLOIYCgZlvLs6WjOoxjUpQP3O8C9IGOT/O
yTBZ6QMKdMT2tP5Z9ouzkBifPj1Vt3HIPpXgadfx8m2bILa51lrSJDpNWI39ujieIc206WSS93cq
Fv0ECcNlTLk04D9v7ly3e8Tfffdm9QZtBQFQAcA6mi8a3nAFEwIqDfQOEcnp99enh9H3gIqFsg/T
TV0gJhA87tqejUb28hTG4gNB/d/XvYRcEtzKBM3KuD4JnuCP54kcxeT9z6WtEYMcIQUYdSWgM1DM
0B+yiVsn7+uqmOGC6qHHzd/A0yqpI9sUBP3Hy6iQ7Cba7yUtZMU8gh/ZP1ZmfJMhEcWmC24zQKN+
dGpyjn06FtUJpZOryJAvAGU0f0sFuLIpK4vesWbfpWc13PJtPBgSm5H9LVTm2g3DpwL8euohnPDR
32CsPviThdBbmwkRQA56/LL5zB9lWS4IQJZ9L4xoNr75J6qEtuXAUk3o3MPg/8oq0kLOwSUpXUC8
00bo1UIlzRH8BV4IqHkL8oPPWXKmMVKV15myxQbcLTIlCH9OzTzUz/dxzSEQWuV6G4KNtEbleNdr
I2QywD7U6swfdqOduT253w1aQDc+aHLbHnnm4ktU2/ZoTn78KqL/X8upAFUECvBmZjct6CX8WTDD
zRkWA1zlzwqpEdnp5ahuWLKI+9pBBtTC5XX1y5dsd1g5iqMiiSu5yjOiK0CpyV99kwS9LCsPfSMa
dyJ1OzFVuO2HtrTc73G6+lc2cSMxdrIBAejSnzk7OGDi2RfLSbBUGoNpoD/nHQ00yWgrGm1RkEZo
aXRlWKKKQ3HBDqd9ex0C+aY3NUDl7VHgfJJv34sx7Kn5MD/MBKQdqObN4FpDqg1y7AMyd6fL03V2
hITnSagbo8wIuqX2/v7xW3PiwkuSn3DDjdxcLubDCBtEJVtXUn1pvoxueOgeoAsrbhr+awaAGqhb
tT0/+PZTDdvX7s10eJpYe7Ro9XdFnSNiZUKqe2K9raRi7PEt1gLLPPC98eXCUuK+RaYwTWzC2Jkv
9X/pL48CX7J9lBGJkIIzzcMJciU9o6jxH3uTly/gS17vmovrT07JKfl4dpGBbm8p7L0eJYWlp6Or
Tkx9B9YoZaP1wKPVyHLxTh/5wUcOGYPVsvipMT/6HhPUpxfmkGcXDFbupPlRNRfysJFW7LgdLgq1
9y77NpkF4cWWDkGH9h6p6PS/7HYHEuo/e9yxE5MdSmwEr9XBuQ7V5VZjHWvfbyp6+1FwSmL1gdqy
YXTiqY54Axa69lVUpEM684bdbwpRlrgEkbPSYWyF/Jvs06YleIlQI0s0oAp+eFQWV0yqT//aWZQv
gaNc6DJnxB10fbNwV4Fi9F2rkzSjFRi1a2a/XsK2I80z+XaE+YVZnVlEpsSJdbykAEIn/qnb+7Jf
I07IPPR/UW2j16xet8KxZpnP2zjJTCVpBfrOrZKNN8QE2cnD//3UM4TLm6bgWetawGD8SGyePH32
LLELOoaI/Ta83YXu6eslhFlV+VasfQLNbToPoT+9JH3PHI1AC0eHEZMt01w7eSdTwxbacgOcMnIl
qoR53la0j5fTYD7lw1HKNARnuODQq+jP1TmZ3kiqQcuab98Pprx9/zTHGqZuLyjDqW4rTF7Op7OJ
AD0ehyZY1C4QmZncZIRZzIBCnEPoJLPTziHxkdn2koC29Q/ZJ5sBJUCscRxXWAAjxfTJEEXV81n+
oDodLecaHK0n52msrJRW51R1s4fS4oHwelOlvC4K+aBlRF0AuvS4WySd7/KuCTCZj/Yor2INI8F2
3fgAg24e8DuAzisCqD2ehDBtCucXHfCfhE55rvbxl9d24Jig9fVHSKnW69gL2l80asQ8E6rPx3Wh
vfMbxkyaORJ0Xo+fQF15kY6Kc0kQ7h9XTVJb9EKAUSV1/HLSeYhNb6/ju/5WBqXgl39Xxc5umJlv
wwiNjke/3GeHSrc2OHG6rc9CGpzHp6xNeqBxoEjc9JVSAmif0c+/IAb1xkU84ZAV1ajz7erpOn34
UF0q06PT1T9AZ2tdy1WL8fK1SgLDN0UU893Zn+3L9ZeDl8wXIK4LfUufAN46djRn1Qm2583grCuC
JVH2nzQ73d7QTxC864HaVWkB71xPVwWom9PsWuqF1gsY1A663X4X+K3+eO+LdVFyXg/EE7TCGfR3
H9OoxEfB8YC/ZRB7ViWLzzLgBBvfvbKDDyGIowO6WY5CYv5gKqkaeeDqrvTWFCEK3qfqsM/bG2pW
Tb/HW0z4SepCJ3pdw4Yj5ujd+JjD3e/4Rw4kGd2NkYpHePYyam4VTOf/gB6bD+BXLTOab1Q0L9zQ
lz2a1XBNB2xCsOU6qAINjNh91FnXLlxExr+R0F13d3nz7DLi8jNGsn9bftYpCsfLjlajw9uz/9Cg
/wbUtdOFsSkfM2XWeHUWIzc5oVu2P+C+vU8iTWDjy3IlYXo/+qINeBs4KHSwnsm5/vR/HM7Pk4gl
WAj8DhARFGWMD4Vz9VHvFzEb+HDKymTDps19FYj3gD5Me+9z9Gi1VmlIwESqrSgnAVstGZqRcqp1
eeDDU3NG9ttjMgFORLel88hvm0R5gRbgasZLS6t0YwP9ZOsP+94gSM9vGxApflp97cT0Z+iNbtfi
bNjEa6hr8+QB3aiqamj1tprW3SzbHDOpzOWAaY+DCl9+EO9AE4NQykBq+DTOgPyCmyTDovj96wrP
MrW4yKIia2di6GdhZ17j77N9A/yAfR1bfI1SrzsQkGdE6A4JjTdPyDnOH1m0cFgBp5tBAfA1CiW+
slzwalS0r5N2lyAGLBnjx6RXWP30313ZVRgdF84YYkpL93zsWPC+DbDmb00PPQNKwn3Te55aQw4s
+HBPFoawtnd/aC+tonB8ON18+CwF7yWjH5otZvkg3P9TQodkHMSPCPMedb9WA3VNgYQDiw7XWCnx
s7PHrOSB4QDoSrM4afpX9B7UeYKCQtQm+48F/Pn3u05bEYLGnRYHVAKUamt1VpZZiNqlzf8EYiRV
tGZkCeBZN+E63HxTmCeYHDWZ8ByLq6fDBPP2RQ0aQCdk5hETShx2kNUmUNoefs0Bgt2WDJxMLRvx
rDK1b7Tpg/kWtSNshumXq+/7lzPVdY/8XEOBb12DWhBQej8e44lZozRKRb9dlCYN43GyPMfG61Pm
yWR/u+lvpgmdz1kdV7gmYCaMSoUrbSy9ljCzSfN6meBEf7aUr5JynyzccmMcQBYhF+yKKFmBas49
i4P7suzoRrVYxgHxYd2/1a7KGrIsRKACwVEkUlRCvgz01zGYXuwKJj8i5Fl1vKMyXchOb9c0PSRy
THbdkEbn6ZdVzYt+O06AjsRb39LUXYnppssFaU2AC0oJaxWHxhh65Y1f2ztUSvEL20CpcFJCZLA2
2ScCDLS0aPtM4hDGmFKTG00XxWOlydzjcn7+fFkl/U/rksb9pZ5oYebeLwiBMRB78lFIFD7FaBeE
8ZK52ED4pV5RtUKRBAwHh3SmqBmZUiV38HKQ+OYyD01j1iknQkfBzKzc9eS0av3nTJ2W2WljCyMq
cL5/yl3gWXLywKH9FNB5u2anG3AQ5ZkXJercr8ecTJkCbBYIFsi+doAlYIqwhiJ0AQzLjft1kBf5
MdmNHh7Dpb9/5AdZtLBsj02qd3h2+AvCAzyElO73m6TyB/+Ok0/LkO4HEPAjeGbVMov6OhCjBDAy
OtIdxCl+/46kSbWxIwXLqubM57oCUFobvCC1e3Obf7cTw92kGKz+0C34SMq3iY9h5tMauhjw+9Cu
7Ovzj9nyu96+UOqg6kpDViWSNSncvYxwaAWAs1kNtaJ5D7XbvqXVAb8NoMq2LDaUqdQ0DsiKYrEA
E/HBqXbDjBprSZ0zESYptC12rfbsVIQg3S05MXNfnXKsc1RvAUYve8NN09SAHOt22GuSnALbS/ef
Vvtq4kA/32t3QNo4riIxD+ng0O/LTGrNJl6uin5elO//I5lwRirLeae3R8mIiUDcGllWl9rqXmiI
VFmWl+njLCI9AsuxGemgjbOaVUfhLfdiUPfdmemqOQUiNi5/HROOi4OniHtMxpjJVHkkJHTPj4ZD
hs9QorZb16bgixMZ1nJTgGeO++UrIzyqXW23C8A2o9PV/YHBpKfh+blO2aSzEMwwRi7h3lEilb69
0kUWvbX3DEEGb5nJh71yyV4FaNcMVWxBZdppFmXYc1kaOI5xeWS1IBMz/FE1U6ptzmRhJHMSHzA1
OYZFt+uHv1VBuVZaYIATxui1KmNf9GJsbu3Tv2Ht2gNk59e7OlL4VrgiXTzAvmbz26uHVV1p6LLi
ysbfya7wNlyJ2ej70wTENBYFyuFAyJFoawbb16tSxxtkl4niHj7OW/FAuJu082YV9I1pyUiqBtVD
cR8KuGeFzGAFmNy21mnLxpvOGLPsuILcfXPKR4qAIec1Pb3Kz+MIFv+50YlMdPHllp8Msm9IGIR3
NxPY1Bt+TE4DJwAF/AIfz880LnuYpSOTIFfn5W4u1CDqc2OZ2s1H6Cl76UcHhDKgq0oSmz+fNfZD
1ZGwD4c3uOivLM4vhxrlNB8VTJBu0kZ/gmOcFpBopwYevXPjpyCn6T/LLFCt3z4XIq/aaQSJk27o
0s1mGsQRMKZsArSywVldvGnmHjIDg4CSBzznaY4x2fuPRSk8Wcil4PjC51TAA7sDzJM4OsprdsIF
QufXxxEEw48MAHwyF30bwKZ9F96t3Q6XfzXHLHQrEwgnpZAWtpmfhrMkpyShvxKkH3bQIAblrYB9
DXdVwXXmablxMxnliwActYz6SV+64G28XKHhcqNEtR9dj1h2bLh0m/bbnYWmJaHWNJBkG1DGCpQ0
lK/8VCd1K6Zp0fnoICNySGjqWIE9K7y5HoFVFVnWV//oIzkgmskyKKigyI+7kRKRwcyEj1cc8bwb
a0srihs00TIz0yHGtT+DpGnhsrjZbvXkXfR5MoOMDHnh7TxCmE1jUo3Pr5X6KlKuNxlfeJTsLy9R
3aeJnQ/LL6tWp1skWTRPNNdx31+rkfHWvIQFZbxP/DB0GHLzHXZs5GxBz9U9oAV2i9nSzMU06ZQp
k1Qe3U17+S0+fkzeYCrxIq1v8rfvbY6ZS0x9vUd6QxKXyPF/E+DRo3u5b/jVmo9E25Qhh/tCYUPw
rma97PPZe4dK71BE9Lj+o8JcxYExt37CS8sdAE4MEJSm2qjslEqoJhAORjA8Y9B2tyty7B66BrHX
nOdfa8dyAq1127U4jSS8mvXWDGPFqDyTy/t5c030fhyHekmQgwCDHlseStaq8fSOw0xZiZ74R0fC
TTnRinvIeVhQ26UblvTnMi2q4lo8lUQKUwlsjlxdpI31bK/C2PUK//qfx9XeXo5XvkNFf1LSxa5q
QOkvB4kMybbpSHCWDn0ZZw+ieIdw109xMJj2rBkgz9PyyEEOGE3Nm7UHIjCT6ymP84NoZpx7o7FV
PoosntSGoDpzmS8MH9rm1PmiEQWqyQ+p5USxLEpJj5COmbXsLvHeZqL57EuJJWli4TT/cKrGjvIl
CFfrz/apVvP9k15+CxXFPNSbnUjIJGU4Woi9W48IRhUPmLOWOtnBspnfiDGFmiO6m60iZIhYznYy
8J4zQ4WdKtmX0Gw+MixfQLMB9M/EGC7D7p+xt/GB7BYAj9KmHIdRssyTmxH7vAk8R0yL5HbZ0Di2
c7tg9tPSIYQ6DG0jJOvCD91CfmXToq7yDIg9VY6q94jvkYAHV2uQMl1ICiglVGyY7zhNGDUZnWZh
9n0GjH+R8S4K5MAsDe7ccNPMQ70wNUdazL6ENc1TN8UkBUKPSg2u27+lq3f/E2YtIpSH7GS0jihw
E6sRXFs2uu9RocsOH3wYT1n2NZhy2N+y4vIoRIVecaElJeru+ovWU4iM54YcSkv07Svsxyt2th3d
0pKEo79kzvBAIEn4/DQb9k3xm9QJ1SN+SpTO+r94MHRqLBDzdBSVTiHLEXBM4udYMjDoVazdZrHC
PamIf5Ldvbzq0E6NtSS98n3PgcOKhXi3de2rquDb9jM0C6A8PjA0XeKtRhj0U6RVl950cc0N19oq
IXi3ZY0tyiBv0z2x9Tt8LHnqLS1+LiUI2+6AyNYGfPWWZeQfJPVTqKFPDRt+qSC5Nx9qHmOCYSol
EtlPjdNSXOvcSljrWGQF1zlC1EhoI5IOo9//KFa0p9cVL9GoKXtNb0phF/DU2SfC6pmearyE1cqN
R554m0RD2htz2OJE1hnZPOT1RTOxhDpp+HQDFqK0CK8wFmv/sOx4wara10ugg1nt93WgnvP0kEH9
+UoUM4giIDQg9CbW3DCKOiTgyLJrmTzJVBkrda/aOqFMtDvg/c1gpEfwAr7Vwl35PHKxdFivI22+
oTcodcpt6AysEfnJgADx+Wy28ymDSezvZkEJxF4UPR0CLi09hZp2J42YbtzH0S96l6Ap6uqWqUaL
1Y6sXaRv6EY0/p6vkpwuLanjy3NiIAeiUHrVdJXOLKKF7A1PHlM/pvtuHJTzRR7tP0S4xcb60Teo
ODnM4CPFkhrPqwulK/QGickU++4btNWcLFX0JyqAcjzgISkAT8APf4U1Gmxs2opYbFwi/LicvNVW
TogE/m6tLNyRcATChS2gKfExWkxEFwGptUh54pKogOnfwVB4CFSjJ7gQPA0paoHXmhj0teEnDxuY
LFdDSaBFt+g4LF320xcNiJtDKb7rGKcH/OCoVZOSQNdYgetgdRqSW/kCAuu7RMX5qGjIMthrmqiF
qgBFm3+y7alD3Klccc5ehvoY3kbZ3Ed18UvgEPk5cbwGO4/6vbF+/0AcvsS67EVHj3op1JJe/gfA
ymLD3TaE/sqwf3z7X+NmsT58qEs77FVpSY8pxDWB1X66iC7IJjYjbvggi26SQzpqzAuiR2qFW+pY
sDPt/Wz2qFszWofo8gTtaaeS1vaFGvDo3Gh2gYkvM9xg6UJqZJLIwXUdc+1bmSMvDTv/t/7tvpRx
Amj1koAyJRJ8Xd5qk/gfsEHRGJm5S4TECsn4Mg2BkUc0S2rmCx45IXaHMOVUeVsVje9QBZKgMAPB
r4e4z+ELcybBP1inIWHWVCI2/rNEwEF50t/dn7kBhqS43aRxAKabWFBikz5kO7n/GOC3h4DeAlbV
stngwr8RaFYmQ/8OK9L2wgc1DenbBs4QCM+8ch/3jAXxfmiSJM7zNakoBO2Ru7qH7tbD/BbpFohd
F97UCyZEhwmoCksu72F+wuRcPRtrK+bSK5ToO43PeAFmycdWjYsNu+lm0JCNp6OTaaCNXxPixrRh
jEVKrrx/9U27Z7SYdh62PIEXhesX+Q4X0Apz7GQI/Og/u44vffsqkM6+6nkuADABMLe3OHE5b5ET
CYNO8MspYNf44qsyg0Ne/mt1Gi8L0KsehX0+uVTEjQTjk2+B5on1OpkPr0viN55PthcrvxAHYpEu
t0t7GxhmNnA9oI76qAcwQ4JAYcE4/spEt3KjXfkRZa1ec+pYU7JeR4IR6FI8kG56Y4IS3HcAcm+/
rW116wmZmrShelIVtMSyaKy74441y7M1hTo1S5YsscUuwKPZAeMqOBLElAPFvBgEXlbcftMYdLcF
zQHYiklOBZfl4P/g+U1dY/mxwaKrbZtbJW/KB9IJwtYcEb2o8Dxa7jmjykyQ7zZxNM3M9ZveRGis
Afo4kf3oGbVdiqY7gOSzcQTOT5eWHGhIi7vpfxwYDQgxFiR82wyqKZ7pzk/aBciqDa6nWIE4gJRU
tz3D5Di7KOmQHyYqF5QikxDlmA9exTo2gLWwtM/EipB0ZwHkLJo58hJgiQ6tHR14Io6EGXfwzN79
61ZF5KeqezYli0bLK34P4tmlAMlU2TR2Ft6FGCJE1ICWbRzWmrcSWn74AQ3UXCm2qXypkLXwreLG
pOg0SOm04lBL96RxBwzWwWoXgI6mxSejSP9MBnsx1zDSO/PH3xfYgZp31HBg9HUFU5sA9rwvVcAr
2kcVWHGP/8aVjW3b/fakJXJHR8pMPJb5Kr9PBvcpqmn0W85MvO9HxaSga9BQY3Iaok/tJ7FbpzGl
Sphi2pdBi8XFuDYM20X1WCUDbh0xh7LZFM9xG0oJCnh5/cBMxVFwJ/FqQEGfrerniTtje6C1A8Sf
CRKwwtwEJ7gUc3yPtfT5g4oEAqbXvhj9gAPjKnIwFSfkaP3bFaYvYwRbe+FEWDRrPCklLLTWAIk2
oaiYpHdtqWKvoczThfhlkeUJ4ALeTX7cedDOquT26B+cMXbh0mO2xyrbznNnG2tRTWD8NSrzKES8
JMq6qrvgnGyBLN1PptUusX2MiIDwqBBpHfDw7NQ6S5sm90ZSk0QhYVK9T9QsWwxjMj9jTmkZGsJn
jCRNccs31cUKnkOt4+jz0ujslg66os41dQeJqa7UsWF6prPVqT7iy/XX9owseUlj9CczJtT1vw04
9mh8xmAUB/BhKc9WspRC4/xduYEgnxG1qVXQHrGRDq3icYi0NR4ZDtplrdn4ghGgAjEjI42QTg+1
QtzzkG+89Ehfgdu3dYuE2lqdVwALZ4zrMj4T2qdv21O97+DlkZ5Snw25aV84enurV+NZpVMIrV6F
oq6EfFArHn3i/GCtSQuNOsQdWXcNVvNfaDxJj0NVlYR/kIqvrPT+rJ1P2HSwpLemAZGyJHLZ2ATe
V9fsTCotqmFb0fvc8Ld65hH+7UsCYXL54b26y2rI3XpeNsyNGqggT9Pr0v+WVeXVpDjw48bTYabV
p/xPS5l1dMe9jb4jEf3RWWJvFYvvztasNhvl5u7VnnRniZHmAwaVxRu+Iunx0Ob5j4Ca+baLokG5
iDCfe1FvzPWiWL6AAGwTNoCkV4HBn/P+9MH4OsMWcLuJcUv9qnbUq4yzgGMvo7nqGhudSTZAgBqK
fDz1NKbB5eiuXbI6L3fyv3RtKzNJxhi9Ex/bRY5P0eSUx0ELCLe6KU9KOE2CG5nDf6laRDL6VJwU
Be4M9KUfIH3WRaD/43Ob/H/322TcXrbczjC8isqzTyl9Wek3nCn1WKZy7UTAnKZY83Jur2U+965u
E2BpXmE45IMoQcJoIjuxyyTpB9oU3drk2YuvsMWx5uF/pPcPS6hcolVs1rgJtkjpHFc8iO4gnGua
77CmOFVBK5fGmsRuGjzmKkoVK1MnrG1vzw4HCDy7Qh6Nw0s7QQGz+3nmql448WfGMTymyqHAvzim
EZNuVZ9e4EwmwWe8zoTF1wTCACH/AVXgnQBZGTMblu4POV3HqRDpPtdmfwc2lNcxOV56KuWEcvZz
Lj0sbS5juBtYGQyB4/5MuYwmd5QgckDHmZkjBEpyojOg/qdklXbWhn5M7ZLepG7htfJ6h/mj8UnS
GZGxX6M18wGXN1IlyCUsEuyI13occgfX0Y+YqAl1D7g7fMK4LrGp1ea6REHei+83Em6cZP8vuuIt
AEbEh0+QoTCu9r5BXlzTJhFu5+AMM9s44qi2eQPqHLrkxxUvGGHcPx5IedXH20l4xRsGxji4vleJ
/0UgIktx2PUn6Jh0uzkJxPwAZ0z46G8V5UIz4SyACViPyiQk6CZtLqOU38msIwZO+Kk3r6WugSoT
SnDAJGnPAMLUqHkgU9dLcjPyH3MSpvpNLAzsZwmdfwcArU6cuJy8m9QSRLrRfUWe3kUwJhVb25He
Q6hXu7+WbZ2JaEbT+4e4a29CCk9hptZ+rjY0Y7fMzdziFVP0ttQK1Ldg8KyZZk0ZUo76sBxbXVPz
qEzyuLS0C+gW3mFWv4LO3CrhKdbgZkF2eAxN9hpWzRv8iyaCWQety+p7U38DMuDtHDRf/FRpk8PN
KWeEZK3olbQgo+tZpyiWHkoASDAE1mOugw6Si1CB92jtXizJ0k4KrhwjMLDGoGQj4w5JCwTUSe1O
+bI931LEHeobx3gadvDlxPYxA3ag9vgY6bzwri37G+Jig06rcV1aGUpSiW/3r8y7S1XKEvh4/Po9
NfwR2J4XLwR0DjQnn399eYVpA3vK9VTjfBartrf6lKD5DEBNxJeC6oc1BBkl4SDmgpkTlBVlam09
tZl21k4iiOYfKcI4EgQnD5q/7B/NJfT3PyCjT73enOq5TaP8Mp0KVs6N7kI/efNwCehC+P55Jb4i
L4a4L/iD6PWxiwXrWv+53ZYOvffP4yroLfTndg4dzZRcOzciopKoK8ScRBQ3GZYSIUFwyT8w4uhS
zkwQEjaJNZeF7tWJFnGJvLHqX9ebv8Eg78UUCnRnTZTDUCQgFgwiyyYl8I/Vhk9dHkgpWMyHi01k
lC1Z66zjcxGs/2ozsZg02o4YuFHW3yApNBGFIc6LEFPP5ovpkhAJDqjQP8T/jkpwxPOah+9K5aA6
RSiOISv+63wqmlcMFpy7gXQyRB6XOV6dYJmMwQUfm2SXUCjBmDrKzkPWN2uutfWbpNI0i/t5sM6Y
0RYJtiCdrCXwY4FCEMxsay7SFi6WOS2Ixoht5O7Mk/Qw0oLKZ22srtTbSUKzkCHYe0ekH/LrLIpK
7uDtLlRbLVL77UDM35GlgRrsCaeq1TGI6YJ8E7ZN01HTUgViG9U3zU3yQYixvY/QSYXvHKds2H7p
wBBszhFAIlofTfvjzT1JzmgvLtXRWl7R1DhTRVE6G909pHN7/c/YltkV/BvXGHYZ87c3ZSljFwIt
uc/TFvmuj8jW5g3nQ2C00qFvBcKoQAZlh4oEMwWvRsBrE3Bm1ADMRbjqo6r87MVOdK/aALUMAx1m
uF5PYWKdH4U3g+08qIgK2yt7FaQNvFCaO1fQ7AFJY63n1lHEkjR0Cj7TcqUiN3vXdmYEqvrYo+y8
e5JBYdvlDTtwxnYynmMalPCr+vOuggXb73uK2utORhdOagSl+UouWoh8ve0tfqVedTVcStsHMJ6H
X+l+tJX49VHCXJrczsdLiZpL9SV6XEVlbB37gBUeGZkIPpcAtg9c2yU9BKLfxAJjSQ5mX4t04EvB
RBsYg8QqfDXkQNKcKGDb8zaeXafukSDRQq6LmgJqwMS8TKst3Ez2iGyGnyNwFmg+wp3wT3FYq6G0
5GG8uPkW8tN2+y8scGMFHLomx0MFqXGnVefwoSf+1NgBW2a/b048B0Cif3Zu4hdDUx8WIkQ4LJpQ
OEKI8I9jqwUU8I3nCMbtE0Pw2xyNZZJ7E4C3LdwmDVyotJ58/bHOiqDezWgqymkz8nSFkILYpOq4
FDjzfD066xFGYFcj7roRnPJsPLH7MSkJXkh8umeJDKMydiMuJ9xzecBHBUc56aXCQxa8IoQrDPHW
okoD02azpeF3Xr+E+auBUeoo6X9rhubuO1U0Aj4p+ki64bAL0TlwjC8D0jE/gb4p7XbLvYKdqU30
mS1WNG/CdEyIEtCM6eGArn8Fg+yGOR8ISqKk7xOknZDBcWSF7CYirBnbk7e9oY9VnAWrGy/pORoN
9+fZkRei3/uaa4eQTjyHNmEuqtETCZwbDI3PNtDf5xG9Um0fQKP1T9Vg6utMEMbTsIrutPCs7Qg6
9t6MEfqOkQ04dDDJHvIXpXphvE5X6vYhcmgA/twYtM/o7a/GL0C+pZ82BIZchhtf0HQJhK2vdrkm
CCPscIG8MwHnEf7rDj1oPWvS1LlwjABAYIJVNxDsSTA628pZZQcix7jTNIs7Ktm4qQpJ41epwVR3
nbcakVyVhNoAHGY3MTPyAThzjl9rcY05KvZkIaD6anH2sek0WSB+KiL4Rey5DzrAaKnff+1KmaVl
JBGEpQW+lrwvYZk07Fr7ngaJ0CPGvShBxQRasqlO2YkUUPiGAFivQIss1KxKhXjK21mAMnDsyjGm
cx8zuMrMqdyQk4ikWwqdeAluUYAik+YPFQIBnxihgIhY7aAf4qTYMFpm9r0YZKcXZXgjYZ0UxMQD
mjsMAeAQVG7SR2Ie5nOj70/vQZ1TBnygNoB0w1JqH2RKJUV9f+fZvhGlnRi254QeUsQYAEGJC9Sh
hl9COx6erVHHE1aTJX6kkot7sGqZxaCHHTym2I/bCrgIJC2nrwXDNmb964ACqjSfAKfG8gWcnyiK
ESYmA29S0coq+kOLJqzC9QZ9QFsaUKFX2bqJnkdsjkT0Uj1KWY8qyJJ4eiJFPHRsCl5Mq60Qm6GJ
7wVKrzri/ijxbmNCSAo+DeLVXXaYP+s5fb5ESnTphweOE4sJoAZHbHA6vKqXwPunQVodoL2lt1rA
sXV4/KMjFDUhxri7Cr114zDPY+VF+xzpSrHeRebLZnrIDeTgVACgpkw71uOahkUuH2/z9158Abuk
Ef86otv4YgvCyGiEVO+F2z0r1tTmYWB6kLOZPq2A4lSBDTJlvI8MUSTM+fbiXBhPiTewCxMiPZLV
vpFqT4qFyvlJdzwLSLlS+eeLbockvhkkqkcE+2NPvS0PFDvg8SQTPGRxw097v2CRpdM3wTXObfzR
q3huWIFC1B9awNTocWTpTuXi7s5810PGxTYFsVgjPWhEiYbjnwv03XFj22ok7t5PIo7rOPiWUq1c
tMw7lH7YS1V3qESS+h2CC3WoHlLPfWVTchEX7r/3XV7yqCDcFJoUhdzatyb8jfQ/oO4B2DWRMLqV
uwU8W39BD1yJF1tYsXW9pjPjNlnFOv154Yl2TuOmbLIYx4UdO1vWed8hvRuDir0pcLg7n1mQ93hK
XIGpmPWZ27CuNSdztr7L+eBXpx2DNm43vns6r8VanXHE1X395A5cyvE+tTfT2jH5lGLO45qXUmPW
t0Ia9FL2aW7YByM5EI7hSvFfzlAKDJO8KGVUZ3WRbMhiss+nuLJ4A8Lb1xqv324YHOlhaD2/AI9j
Ec9ADKShZecm624c9zwa8MG/iLZo1VvAgbDrbq475fPuVdGNzgAV0M67OMv6MLA8epdRXWj49B63
RkMrS3q5M0KMAt6XOqmN6tcQFaKRsOtZZqD6DtZFKfqUo/nvJw4VOZyD28QC/8yCuWKjkO6QLWR2
riYcXyktXb0jCxeQw/7GJkTuDbQo7878uCLYuTJ16D/LFTF7mDn71Ws2D5DZhsFL5Z9kwhfGBQit
PIT6Fqj9e/yN5//arBjAgS5JCnvAaaT6pl0+kA/aeGzaZKezgn1O6RMl18e2vAuFYHP4gIDq2oXd
LFuNJDQAIisiI5A/yZ2Oes4aMXiJ5a0RZdquFKGquBS6974NiQ2RdsxY+xPTBXfUcKUGTdtF5zV7
U1OKhDKOUDDwSFWlWOTsdU/5fxr3AEMxMmc4WF9fQKrNapm0AXgcE37ojv4J+tbj6oaLQqmwR7pR
Nf+pdMWX0LjNJrgtsR8esYnhd7GgCArND3ljo65CY6zVn9y6sdyhu5nI5Bw5XyythKPCqZfXNGTD
ZLvvrjaaTeSpXtptqMfjT9k1DXiJ0UKMikwRhe9CFdhPtjSbXcor6D3B+xAF/12B/ziPF5AMpSqp
arF0Lk6iAA8HTcY8XV1eCty5I/yjTSfluiPjhYxf54OxR5R0X3komH/kGrUqMkwoVCfpJUMI8h0A
1yRGSNn07j9tWsa9ooM6W27X/Y0t50xPDGZe2oALyimf3ZaWYHxFMPFx1GjkBZDcwnjcrzRYEmUV
e43qJYwT5wmmlh6GBvRk+fCN0Abg6PDGL4YAJEeQJwIjaD6qtIFYA/Vv66kSb5fU1tAeLtawynIQ
OYiowGErADVMyLqJHcP4Wrne0JqkR7eEwTzcMuKLkbMCbIMLxbW2Ujr0QWkfiDQFqUCqLfmdgrDA
d+OkioxlbDRKIgxWt+7wAtgjj42SCrNMim3znUZoK975eLzag43SarlLHrGDhwicVZk04kOcmyU+
/PBzg2iW1b8vuJGjfBokVRsEw5sZhIUyPvJ5arJr81yRkgYqTFVObxs2uHY/kNJdtGNw5mbcQpSq
Wzd3iiVWdhBlyJQA8obUavXHQHPTf/GajbEixbth+qwmzSqieh+T3VMWTmRi9FaFbogcWJa03OMN
O6gvQC/kmKhcswE0JsAHeVeV0Uio/oJnWLac0HAO3sIPz8xpoAuNUWse8VvbsI+K65PpZNFjgsJY
1vnz5E8GZZq0zjtTocMFuV8dXxGjEOzxNmM8TBDl+X+x2gQS701maAjYxmuqXyLgYkCWudk12y1O
qkHOu3O5B3ZYF+ayLx4pBrqzb9TwCBJksQAE4M8EKYkgRwug3CUTe1+/w/k4XYcXsLQ6pFWXJzcb
clw1Q4FC+3sQwv5c3lNsEA/YKiTWm2AkbrdB+ZeuNSVDzq6QSQigfcn3SRlgN01ieUjbmdREoNlJ
qXBQT4R752Eh/EadKk+0GtyeQH1+ZZDhjiWI1ytJedMgCFD6xBrmOtHPDrhn/kb5MJiX33xX2dR7
qOUtBU2ZPSTwjQJsnvy+hI/ZK/6wXU3HT70ULlByQIlpwQ2zXwv0fxQ9ijqfwgv1Bx6RSH70I8NM
qs+F6iAPvAAkyilPOyUlw/4xmceQX4IyyYvLyxuJVz4OQW3to0ZLUj9l8Z78BaDh6cjfEazZ4ieQ
KadEDM6Vvi6eR+09Yjpp3o8h550pU8PP9fchDO4eRj7mfxyYd5FyOECJADyRkkdIO5FI0uulVAWK
hUyJbGvxwZMNnZ1GA83F1W8m+ceMlx1GR+qtmg3dDGpdCOWt0XmiXi1AlFF0oneucUfSphNQOFER
rjA0wRMJxIR3kKLB0bF8JYY1hjO8ItVl09+oaNnURoYkTziVspks/EByXkMvvyvJD3M0JkM3/0E9
q2Sl8YcqQTR0n0qKKUjNlW9JCZsUOtalTcXFNRyhkQzHgS0rp/dzjNdI3Ongha64BLKekT5Cx3lr
I81tSbDtBMulzRb7U4tGHGRM4EQnT1gwIuqW93iN3QrUH544w8CG1XhYS7F7r0AsFZxzOV1zk24N
0tZN/r5vlys6S44xmOoxZB3XUyobOTzB8cKr9LZNVcci8Yt5Q8oC5+vcslReTtwWKd82T0WabPDZ
kMaTSi7kRPwxoUiproRsHA923pJK7ugw5r7NJghC2HPMv3ojaYwL0Dl6sth/e2SePza0atAfYJ+U
lxO2DqVD9erRk9m6kTnSJGATTvQfDD3F/LN3dpi1PDhOafXecJimp37GHtlNQQ3EjnY4Bq8UOzsj
qo9wKc/hGIJ+cuV/kwSbsZaqXXu66FV6Dy2QX52+zn5Gc6TaBpXe6F09BPqCPAERY+zYYfrTLdt/
Cgwo5bS9z5hzQxWGtSb7S+gEc8VLslQmBhNVedoRH5JdjXqGwX9d1y2kmqBm8zgrNVYpuoLVEdcF
EF6Df5azWUpVJRXaJt4F/RiFHpQBPVRZIsK7mdaz7wLeH8kDpplF3ATssEf6umdTz3gQC1OHqGe7
iKILAwz8yHAirOO8mpfw9TyQfZ3VU08aGXynN3OkV+cnUSjq4SRXLH0akNWejdOkEacTfOmjN5+K
R+8Uo0jJcXWQQXhzGvWnmPoEctlsyX7blgbX6DW3y9tV3DVCVlH3ZE+YtTYwmr5r26Qqvd//s5wk
OfRZ/qIOX+C8LbyB+eQs9AxMtOgYj6sB/5IbZgDbxdcfbC1KoNeWVPgorBFJFb39DtdXcW+0XFBU
+QdNQC37T8jmxt981TF8euRggCyzjTfpwfMb3Y1U3l475DR2/CWDtbiNlsV9HgM7LlapcNSgT8xw
E6Qp/DtxLIW29Brh2GSuKG5PIEsuMP9Quay0DWq/pu38tMBF38kufrAEfWlgxse2Z7+SFh+UpJaJ
hQ4tRL/l2qEvW39kUCO0PYI3ebbJZvoBX86z2xFVPmE9tU2m+Nif90wWhOFfESAdd3HNFzG6IN6A
GpQOVIf4EapYq1x0Jd2zH7EIAL+XlsirTdPt8efti8YoIBy+Y6KTWc5zChWu5EyKM+obi0x88kxS
K6pj4AR7gDtvHmtfp/HgqlqDfi8ggY7A4N8wKLy1cZPly1I+mdGrBGHxqOWiqXK/HgPR1GRdhtUr
DiLbtjf+hAKlSVFysQ2Ov2ZN+8r75WwsKS8dvcjC7zDo9xxsTArlIPZfcciqmENUrzppsV9hePCw
QhC5/oGP0xpPcrNig6acMV6H8+dx2CwmhqN74/TaFzqU4rfQfyXUF+6lvghvHpUJ2qRRLCioFqu3
GUtaLSULqeXyVpcN/YResi1D5cPSZuyWikPPu8A9JEX3O9+PhY9CF4sqPmpOwqTNWVQa/t77E4n+
BeUqU7K3E96f96hUpExmdNMSMxldWEkhBFdHZlL/fAYh+NlFOdVXZH4j06HJIRXplVcOH8lNtyYu
e62MekN2KSFfKstmErtRKWxuWdR3Yw/fEggIsvho1ZWRftPt8iAPYlGZzvpGvwVa/wreSNGA+x5f
v2HW/yAiaWIty8NPrGXBZy5OHbmOdpNgcGZ6IHkjCAuS3M9LLSnGxdTL/UObAWLgTpycadTb3fWT
6M7FK22XD8Fk2s7xxs3tpf80d2+vnF+jg6Oi2Y96CRWe0uStTQOOv+6Pp3CXoXvaJQzAFeMMyjyt
uwPNUIfO9C5ps+H43b71Ex1oeZuu7bSWQdOKmHgLSQkIZ9VmdifoSAd4sXNXHvlTVKrFwRrdrAJU
8zXm3yJgIprPBkEQruyqEs/gBFS4za1v5EtyG2B7BT2Ec9fNCRcovb43YdY6jD6JOjdWAdf2fm0/
aqXRG5+5f/VfpMr+TzlYQUqswitp+UvJO5Ns8dYe1IxSqIsUP1gWmraPr1mGubc/zWlw2vdaLJL9
XRblgun6RMFmTFjkMpwL6ulyTd2mFjnMvx477iTz3RWI0+rlCJK4N1gAyjfACA6BD28ZURuauIQu
hbFDaLMfqjho1WDWmOAPDN4FZxZSHzG/ulfN6DJyq1C5j8lOrrsyEemopygTw59c7jH0I9xPXqZ1
ftoeJISKffVHi7yaj2CDn+Z2bjWx5gIH/GY3nijXfE3hos5r5kZN+N0KHu0p4OP+OD52QtZ1/5SP
qKsl2BNYix705CXO8XoBj72vfWQe8yuoptqIaFQhK0j0lJKZLCdQ7NFKDn88WJhKFU2eQYlYETGj
sZsZldWAOb/oyEXVoF4R7L9+pgCHHoI1pO/VqMAZWmt0f21bWOPheP1bn4UUoH8NLAbGfV15hnUt
dNL7D7dFw/u9JEXscp3+ZqB/BQSzeMN4PqhLKiJQoMTOQ/wY78A+Zn/UWTS9KGoKSaRHNK2715zs
Y+RZJ2Otl2VldPguJ2L1JwUZ+uXJycLRXupTu7EhsH4DG+SFFGbrVVjAJMfyn1SPV8v1Bqa1nGah
s82GU9fO5XC01CNq4zbGsYq4cAtm8RimVJ/01oAfiSERHUP6lBc7E4ef+SL+Ug2UX9edqqc8D43t
EOOr9DmX7JxUN0K+k217B9dxErNrZIh+Pwvhnbxmv42apDWDRVIZ5GOk6xgC63st7YdyDkoBnKBF
3o8lvLiLDq4XnwFWcVIy73omM9vwsnQ7TXvfdVN8+bJ4BWd4gcJ78Grn9SAQ49Ft9xWtpqATwu6u
U4KbySATAeGBebXpmUrTboi+2dn0eS6gspUYQGzcShYaWrBAg6K1BscdVj+Z3zBdAcMjuj73l+Sa
PK8hE1Jo8DRx3yZPXtE9m5yBE0EciDEcXKYP1ZUVVFyqBJ0lzMsuVfKFS1Qkj1AIlKnCpvhJ5PRW
hc/CjgeoQb4GIs4eWnP/7iX3ET9GEc1WeRIEi8N5nn6tf1Rn9jD3I/Cu6ynscVMZYr9ivI2YRiM2
/9TX/rQeIUlmhdn1yPhfOGQXRVrD/6Dqsh/JjrwZVBpummI1bChROmCfjkFvxByl8LOO72K0CKaj
bi17xAksD5WYW94EOq2RuIwsv7fWvyXChnRf07IPopPArFbPRHLq0iaVSshbFmVuipFq4CTDreOr
yXwdB/Oggb9w0cf7HZad/RiRi68fdkMU4+g+Bc35eX19cTYkaOUJ7tDRyhkfzrCsCI2clHvhu9p8
IdIVoly695aLu1oXnBIKoiWFCVHUGp5HUs9lVWkYKrtIdOUEmS7L02iOrQabWSSSRdLZR3UuT6ym
ZYHaEw/06TbRjIffnYckrgZuUqad1tGWb37CRENHmVSJD4zKNOQ+w8iU6hST8eEP3bVVPD0qd8ck
iYEHQYHIqVzaf2GmOaUBF6xfoXP2mOnAbMkSe4Q9EQXfAn3HPKGeUPwEHz7kVBJMiGSai06ptMyn
IK8vIpBtOzulilqE6MBuKVfs6IPWmXkUr2UQIY+BXa3rNagNw10oqGlzhEgDlewswSzSmLlej4u6
4WTg+ggk5NTC+Jnh4aj8yDSNgBqVvECCkeQAytYQTdqq3ZJoCUfavCVDrSvKz9Vm8d4H+HAKjX3N
EsApgkONXG4yTvlKYOQRFvW1woRjCRw7heCa2F4zwhg36wM2uqbgd4jkpq+uuJRPwdAGRSeBqqvR
WpjKutdYJ+ubWktNiRciCoDciMjiV9iBVwY7XSXuyDLS8NX34GXdeXVLpMMCrvlK800nI3xSDpb1
k6K0pFfLe6dynsWenP7VlG3Fu744Y4Pk28J6whOlRzg88LqIZQY9BKeJsDQsoly+v9xKnBfozOq2
Jp4rvaKyZ+n2fvxxw3Css5raj2ihNZGFC23HGihHEGNBt0fNVeNOBWnte3ywksnXCljjvEdIjEJ9
K3YHyo38Neem5CDvAvFX+u5bz51GrAPHrBHlHrBuiSKZmVuWSHygzrFBMWKxEJVLp2LGDR0PQ8TL
avuf8Q6ozQ/kP7tAyBJ1SBpBan39YeawIV1rYU1mRDhmtbijbq+mqnUDSWcMep9D4kaTrWcVwsjN
y5vCfJAF+1A/zrNzZbX7T5GCNs5MFtUdvcEUrHgThLKImgQt01oeIvh4O4TG82bU3Fd2zzNx3hDY
Dhp+U3PMJZz5qVU1zCfp1HC0iJmEU+kQ4tfHfNkV6/GDVEa01d2WNLcnKQm5UwK2GT+GIWKxWPmn
PcEqLAX+TuXnwk7Eaol5clBJ7EctvpbV5su7rULfkfdbhMuy9vhU0MvKpos1CBbrunqYZx6MMvnv
iWFv9z+f/mjFlz/oXunb58Z050NSbreGyvyZgDRuMvsl6t468m5IfOfesIHQvL/kme79aT4vri2l
Lc2BjDPb+e5sYW9o3mu6zLnGI9Qnu+u/M4zu3BYF5JCdb7tjX1SD9rU0LKT+cJ8rWReZlnb8W7gq
IkzXnAnh03vqcxfHmC2HwL8mQwkgoGiSQSX4ytkEdMYJrS8x7sBdots+rLn06hsBDmINfV6zi+1i
cnZdJch2Z4E/71z33aW1TGJZ7Bt5TdkG6TkxXfi2i2oErvfpYvhr5Ytea9ibA3OD9RIFfNUs1DQp
WKBPLdLsesG65XPfo6rwJuWhLELiTjThqxyqhN7PbW3TqSp2qUk+RVCZy1O2j3+RuznSQhqW+ccf
uHn+nhBAn5Za2iNPbqrqKXGm+9LZW1HHxvmv72nUxpCHKRu8CIvVwFuayFe6kgO/WN/gdHMhpJcB
HIpccxlY4vX78BHY1zmhX31fZ3QJtiOL0k+3nNBfAQA/u7+WUaW9uXGXmTX4I6uj3NF/6jgOegSk
cJJPN3lnSe0vv7CqR7PgoNXb/YJ+qMbH43HmyBe4xHzC3+kAbuVznyrcgMbMxbUK9idJ5XTpBLY9
enx+n6PYG1cxjhy5a+z9+nBH6dBxdUwS0leY4Dxhybk6RrvdbFs8wbALoDjMr7UQzLSPaa1Nl4yE
SJZSg7ERZquSdBPATAhjK3sNyahUm14odtC4mlGGOmvVRh94TfkKBGyCO+OOn2Gdw2iU6FUdE4GN
DrU8E5nGBjjWWUSoxwSownvRk9nagAnxe5LMSkG/qCLDAE9WtoVkdrqUALW+3RMg0vMwB5amGqpt
SaYaH0tPjsRY5I1l5zGPwVx8P7Fhzc7JmrbutmUkD1KCMvjCUjPQbCxKwIrBO7bi1Bg9qf+xeL1z
0dUoBFy1jv5KN4YazGBbY6IDn+PqSkPtt04CNN+V+/f77ivDnBZFv6F9i79gQpd0zvCGX/u+RKof
fcefZSItoQkwfcnbL7w10tqIldv9dTUuvsYzgyobBPPb1jfEzvvY07w8hAgambUxaiF9HuUDDvgs
lyP7K78JO3ravBAQzcC0ifksiSQupegyG/UBSPtAyMqYZ2omlp26DvexMG4vClKvWcaB99eN+4Gj
R8KnnvM0/dTSXqndy//TtMFa+MJthsDaAVeyrTiCm38JMZeLuza07KlfLxzrcseiqE3HXoCNL8z4
HG/gM1hDkVwKp55Z+HGWIuZrGTv7aeAxXG0V/+h3tX6sLW0hjKZmC4Km79YKvvHfkpVnWMI1Q2/6
oxJTMMYOU/7NXVnQQ4A/oaDKeHs7v54Xwv7Hqu/k5IgCE4C5Rk3k2sOZ39/DsnrWN+GD7vr/omey
B3HT/bffzF8EMXQpyvWpQRVelW/zHC7bFt7TEUUkLlFX4Gsfq+3RgRrERmMXKZjykbh/XdcXJFUS
FzfWRmn3MWedeCmtiHS01IzmPWrDuacOLFm8n7GgX0VTlVbdY/yCf34YZc6mLC5SLoRJXsmEyJux
nHwAsg/HPKG2IAyi1N2vTA+98xFXWEASvQ2rG6iBNuj6gvbrrDA1Tl+eq3O0CKsUl/RDLyIjxCoX
J1jqebwirC/U7niIwfr5PgODDggP7+GjCZtJaXBsQay1LGjt+x3KQboZS30qPaUPkJBDhjXdHZYe
V4j6kukSfXsqwgnXilCRiajAdXS+41EAWMKSoGhovH+srt4MkFZZRhDnLC7FXbz0yJKIVgMF9GEH
w4z8eNCDlQy5pwg+CoFk+4EMbeT9JOHkFzv2IT0tyUoY+gY47R3XqwgON5rwcMiczOy7vSEkqDrF
o3iIEeFXAQip5YAr2falv1a93D+5sdbvjt6XMlj9Oc/zb5XDsOpJ1D1Ehw79ir/z2cCu9kTiiJ1n
QR7FbcUUBK4zdO0jSVK3FRmx1e9AKCZWwKXQ3Q95/UQgcYdgcx/PFGAXKq/9QvukuFYp0coFlC/V
Gv7fn95szoo0eRCg9M7Xbq52MztV0jlifVPKelUSvfgB5z8XAMqnTJK/DvFb72yfc4n4azZua7lX
UFY0gveA9+ciphOIurHqhtSgRSf1XadvG3WFmSSBoGCL2ORT8tyZewpWR8lqQh0tgaw7ING5lZDA
+j93E5O+v3lY6QXxvgXR9Et6J7k93ONbmqeCJ5UBuvGMqesO4BpHZ3b1G8Qts0NPvg3+t9y0E+JS
iO2ZKXQyueNY2tVbU4uYLHN+xN4u+ZZkquKN1Lpk2+POy+/T7yqw+gLXcJIcUBOnjbaruBXav5gW
aAYMiWb4Je54+z7sLvv67EhPLI/K0LArRFPGimfHwuOGReb619BiZeP1SerdJ0iyC6GeMU2IhdsR
igAoCXrGYaoe/UzTnREQhfE1CttHeqYEY1Q1G0YUMvzJA8HMBbRH7mZcexe8jcZKc5yotfG+kgrF
eYl4wN/T/PTGMFZlCJCXzpDMkM8X0JZ28ef0kBlaKvPMaYra5lVdyknX4lTGa+NJ1deQRzf2gS4n
vc5+NXoXZlE37Q0ni2pUz/021ukvL/PQsuryxenqgRi5LIHuFV8DPqTjuESCKznEKbiIWAbi314G
+wReIDY8+ndRrBAccKbgOh/OIT9Kh8wFpyUVn7mE1v0fPXS57Op6oqcIM3p+wvMrtedYmnvRd45/
tAb9IZjSMoFTEGYi4Al8lZARaLrdtP/b3ocCZ+35praMWyZllyPdVdxrQRZ768Kl61yHkuS5pgvO
6PIC979ZdcziaaMm87vFrCJymGrhlOlf+xwgp0AmbnLHDByg1ZxYtQw6cocZFtJKC+OsIzgkM2lH
6RmKbmNAy/iWV7UdSQxBQiD48WONsNxtIu30CLjy54mwcIat2vVLkP8R2AW+7+thja0+Ct1G+CyI
lnv6EMaA5gmQzfGSa8S+o232whKIYvgs2gEjImi8wJ/bcGf3jIJQ73orxTgzM3+4083upPRirS4I
ZF0Vgy9vuS89bkl2t2qXXPoW5OFPtVIXUNtNgQJtkX6vkGzklJvjM4Vghncwh/Z6ngFTGUQfT9nq
rjUx7szTeytz++J+SgjIv7nu44K4Q17wtMoJveewWgQYWmVNtgGKueejoNmmTDKFk2EyQwSnX2C1
FYJ6oJqp6mibwFcwI0bFPMhR+Cq8geS29eVlcq+Ef/jNbsj6iCH+Odp9SpulUMAC54MJffWljjCN
b5T2KMQsJvxrY/2VBxhbpjCc5ERU02OmVWId1suUcuQ2UjN4Y+YmArvH3n7QE1YcpKf1kzPnvPly
EVwAXevLEnT+SvwSEDnlilnKE4Vwz4U4rNZQCv4EoOSuPxZKRULUydL+TY0rK1/Yf9ADkslzijNV
LEKAnjuV3iZCqxPlpA+ImYTViEP3j3uZrYaa4/Pyrh9YpaUrc1VoEZIiHXu9VfuOCmEa2mebz6j7
ndKVdUx3mJOUE4OjYcEUHce/K7pHpN5WTQAzuNZYlZwfWszLEPxJjXFmL5cBHyorADi1H9e8wsCX
cXUH5h5yOVeXXGH43dfsf6UqhyOkxQPjhrlqKTGAeuzf0KtgqTjdQq5HGwa+dmd7V4QPEOrJ/4PB
1DKPc++u7CLepyC/KUdKsdezs+wgnYJtkxPJDYcTGyqn2Nqnyt1QY5NI25QVMwNNDMHfmWlH2wKM
LsOnImAfWP38+0LpyIr+R4c4HUuZZUFiwexm4tJFmtBnaznrJb0x0TMtgJ+MQTseKgFNpkv34+VI
o3A0oaYcbk5VS3KX19YQh3Y9MkdL0PeHYND22QNIjU8C3kB9YnF0xkhsK7TtH8m1JYDeptaiXrr9
Af6y0CDm/IpXPahS0W7dAL1dju6ahkZEVd/QSUg0LtZTgOcIbotPpo3cjCVHf6rryTkrLMhUmfX1
FYszCCgUWjzbvq8dqvwUUsofqlwtMWr8WSyVndDN+6nNobi8DZdrdSrdgFIwUyQ64rCJpfpe2wDi
kBzCiSU262fscJw9QPdUWqPijUer2LSzay0c4obLfRhstuqfLSSE96IUoxz6IeSt7y292lJV1Ol6
APj9FhmuouCvMeErmSILYjIJWsnv6BQsNDlCAro4hIjsc5TV5DMV4syGoninPpzM4srw+TU6mRqp
KfxQB4p6EEw2QTe1GayTm8HPPHEfIBShQ2c4ayqBbo5f1z9zbnePToOYG/ghOcuS98c4RcuUEkKY
gsZ4Dv2uzbNjHnhUxMZ4Y6Fn00Iz9HSeAOhZvruuCQJXm8k0s7w54z9einougIj7lHB0m6gnzVej
9a5df7Ldo3Qq+0TgbAPrJ9wWk3q/RiOWdotFLogeMqEPmHEpEqpJIIWPp8nvcD8E6dHCZ+G7RKov
QT4EX468ykDyihxrQgQMzXWblBtlMeKquZs2czrMeGqX/ann0z0aUiGmQg9YXp5+L9qKzH35VCUk
O8FdtKBH+wfQUSObZqP8IFx3CSN5yBbIaJBMf9sCIQ1IgjMhbTHqyFsWe4Ri5MF7F8YQNXlmqxje
1APS/qKWVQESWMLdkiL0mH24MbdTLRGQDXb5w867GZhYYmdA3W2YN+MJmDHhHQgwPLxA19/zEW+d
9B8GHqeLimuETIpunVjLMxogPoY6wQ6q9Y46jK+AjfYYRDcLOzLxogtYII8jwWBgceSD3uaIF5kk
ZNDhMDlztFd1boP8TBgYBfTNZ+9tt5qkRn2plogJcb1R1kVOfefcaWv/pqFpYwIGjtSDwMivwWuw
kT6XWllXwotjQj889nenuY5CK0pKcHRS8ZcoBwanGnxhPzDspnM6/RuIDpJjmLhPConid29kcfjA
qoY30l8UdmKlBFaE9zj9FhxiNSgS4nvkBQrE0d2wMA10lQEm2KkPVVM8O/nz0HRJa/v97u7JLS48
Gzmh43lyNdSKJ2jJNnPw+Ej0iTK/Cot7g+wIMTwjoP8yho4d0w+Z0mOdS9O+QtIhPSAmll1dV6bP
1H7r9wGSJlhJsA8+85Vt1kp1TgyAw7UeiG4JZc1sG8YU+BEVR1q17XElbSaHh+RAjkOs/FUShf5K
aECIFdBG8IG/Y1gSLUftIRayjeUoQLQrcsLx0aq0KoJe5q4JeCfFC6eT59nb1zBEdj0CrvBqu8v3
flZxZfhImmdeV2qxlgZXEAtsO39W/FYI6HeU+PrU6vjnxITvM7sCIpf6NcGa/tLmM2BLF4QBg77f
izL4zIbrISYOI0WCFeaGgVeEBX+lGlWDX2iTHrKkZvGHCkXQlC5fD1JdAj5cgHSkaF64Dr1AXrcP
ZsvJw4+iaGW4Iuat3lE2iPDHS9RIa6aABjWvlroiTU92OWrSNeTPlq/ZhpNnKHNN19wGKPO5RfFy
JmtZaz8UAC/69gbo3Gm9dUC1k6yjDdR5WKYbUgID4qilf5Ryj6l2BMBw7g493VSlwtPdr3+avjgi
1RectxTvEZqBpMtqsewZjGDA+YUrH4IYvSRwxjuo9Cjqu2nQoLvAN4VHbtmJpHwrdYESH4FDsL2X
2M/YvsnqX3ZPrQozDC4jif2jMxWAA3K8y62sVqIozsuX5KZzS+qAdvXnvgfCxWe8ervj/nG7YC25
Q/ihMcqovwEXDVpOHLhmV+EvTnrB+OIgG74vbv5zaEluwhRsrFnk6mpd1V64OCGMdrIIowO4e9x7
NBiQD0fA4z1d1Zip2i823Q2efxA4ucP/3U+mQBnEhaB/2+8izgS0P2PbjdG26eA8OmOpeffS3rfC
ffZNQ9xJvtgkaFSk+Vmup4rckp9ebrmdm0yq2kjtkejAp9dVKwH/7Nm+F0F+CdeEKo6sCRktCe3y
o+JSLbSdd/T/6EIdTro7meTb1l4/CI6ijJTVbDob6/DxA3ZnUZm2XOE6a2Hj9z30jfsmtHKdxZzB
X0TOF07QJ1cksW1Pcs6ovcsak6jAx2czbBi3aGssBzCyabxFEh6tQ+bMSSDaCZdVDww1E5EuVO+P
zo28gwbPvqUX5YwLTsMAm3j1gnjMpdkOdWgt3ET3t1VTENVeM58KrH8VXzELe1CqZqt8dzDn9mhV
kekEa+hYtDpWV6uHX6djYCkWXt6E1fZTL1LXPni1mOZDV5Ek8CNsExlguGpywTTo3uq80X2FkR3R
0WC8BxEEiX2SBRjtQcGMpS5Kg4a58V4PCBFTEG7IwvZDW5W0Wz5IaFNHjNnkgB+KCcPnZ5+B1otI
jZDacPrW9aOT9FxZsAwmqcMg7s6mTLHXyt8YDjEYU2jf8shlKibDg5+RThB8tmNL+S44pflgHz8Z
1GFvHuACLb+RnvDSR2El1R3m9F7biM+PpBu/LyMRYV6fGUql8Pu1J+PITzdYVHpL7Rie8+4ubNUT
wLg4/399qPQZtr6MZqPQpDO+91HwnuZhl9eKgQEZjveS2C0Vvg6br6ut7tTtMcxz5GF/2sUxS59K
zjyYuGYduT3ozdffP/Cv67K52rw5IrvbJzLHW7Prb1MfHaybhz+bTbjQimH0rBH/IZbhfRkckSMJ
wipmMr+iO+GGxVAmKCpi8dptkHeu8S87fibABc9h3ysmYOlexwXRlGYhfpcjeKhza59jVfC3/Gvi
DiVRRHKbcrhA8eya7XsPUMHuCsLsANU0M56VVwBoG9JBFGA4BTl7X+Wre71LITh4vc8n5Vmdy2kb
M3pz0yReRZMea9Rp3LD4ysvuvutPSKM+rszSQ4IZgf5mJ8eqPj/hjA08vvp00u5IcGgh4AtI/cyM
d93MWxJqKT6BcFgibQmW53tYIZbOeFdEgaRF8pANKAdkdoHXE6Lmytm2DMRXVsKPgO+/cC7Yz6he
wrnbdUlKwY/6h5klblKOhO8rDVK3WMUezqQD/2reWK318m760uYS9xX7D01rBqzMGqeYkICgnxZO
A54galWMF/jXevGRhBxpNJnKOpW/J1Ulxaht0gANSDzCYw1HSiaG6dccCqEVxm7fKMCZ1x7fguoU
CNbJDwsVX3GwJI/mqnFB3ziGvRa8RenSJi9RzkYJb9/8f5jl1cL33b83QHqcV0M4XWQ/2RwbN3rO
TqVmUz9K/IBa2N3t6rq1s/dVYOdb7RS057Ib3xIFjvM9Qu3LVZ2EuToIVw2PYP/FFhjdaaOtJLNy
7YoTgM0A7ZBKqK7ViPDmoR8wJedJ4AJgfbRrUpdR3SvVvyLVAs4dRCRD+5EbsI+U40O8xY2MyDql
1zApLZi2cupk7pAylwUfM5Qj3ttCzdlZKv/0vJGR22AOL9PnnY7kX4oXFSC52qn2z/B+5YrzdAKG
CK94ghvT2RfbwbdYzJXq4ye0HB7dWEzlEwvffzCsFpgSzCuVAB4SolnBoJDjOqDLjiQCj9izY+vI
TbfobbUvV6hq1FoDk8iyNHvygSVmL+rBz67PU6ellqPjc5jWFyUT0OyH5Zp2lWaZwoc5uo6ZNxhx
a6Mbe4+BjUe/lpyfoOzfin+M4JbCpZ5/tASDUNuGpSjq4M/3bKt4+QvfRzfxSamaDC49tT7IZqFW
bMU/i4+45g4QzQwh48gh5e7YawgrZa1SpHBnOHhZja4wIJSxwQcN2j53bqWC5uGhjQiPXHKr0m3r
1F9T47U0U1nQqpdsBCqUFb0nIxL1k6s8I3cf7skZvrEAF41qMdZtdfjktqyqiqey7R9XrdZBm78A
mGv7qAIrYYHS4hXDZ2Gu4S52liHjbSuetFxITUO5UJU11J6+nwgM8tSbjLDy4qOp+y3+Y8h+S/h1
h4RDLH63yl4ZE1jTVnlzXGJobNEHTDHnf6RFcyqLXjUXTR/NrO+AgzUFqDulLJXRRu46eou2MQZF
VbRNNnMKLccz24xLbjdBZ+RxQXf6P4v6IgFbwdb4AAuWYsPwmsnuISGcAMnwDpft2ApSvUQxafCo
ky9iCUFnf/k5a+tkToIrv/wRtzoaTtivBvWDawoXg5GIp8hVkAcsSSFimFKyN4wEkYIzi9zmf/1b
VFhfQky1BZojGzNybjxjekQ6Ul3m063EuR0jM/yiPNK0Ncafkstg0HrOkFh9YKH7pXIl2DQWHBfj
8scWGjRPz9i9Ap7iDoTjQ8J5CiOyYKFEdd2sao/T/IhluziD80i1j1RB7Ag586O9Roeiszfmt6Ln
4eIseZZAgC2Ia14zz0tJsyJTmLiUGFeGZvcnHXrH7wYJCjyoOXt7V5lux6C107Aa4Tu+oSuO0vT5
mJJF4oQnBlx1talgiQflkCIGZMm0x6lEb5GPk6bM/Gf8GdzItzuMAzYnpc7POk0lxsRQXuREQDQ+
8JLXB9MjfcwMfhA5g1/IUJWrqROWn3QYFiOWmO/QnbOglK1BnbGNUFtYRmKbQM1FV61RwJ0Za0o4
JStcvmpJKpU70mG7tOjwTV7smhawgw6R6SwaUJ9bmXQ82bd/sXluV017BepJxN5Qd187KQa/+1Rt
+yyzA/22OmXdQSG8j+kcGH0Ksx8HByAcwgWKD0cfGIJKV1D2fdEb70Lxd9alb3Bze+NZmnu5ktxS
o6ym3/CbvvYS12detS6D3x3CIhExGNA1AmVLB8SUyiif2Lpio//gOEfgHmL5neFqEwwgoFksJVtr
/yYYFe9WQe2Tn+3c9F28I6NJ9fFx19rCykKtzwvh6QvvOusjhKwbuDP6H74WKoKoXg7uHqdrEErz
rR5cuRWq/GQlWZN1QIbuN5dXiyieYQsLmeFQnfEkLxA+/MAwi8khZDdCzdGNvdwXZ8qbOtpunYT6
9AD2mRyIYzg7a/4rNmhE+983kx/xcIGdK6deH7+qqp1v3w5EXa9Hd918RGAPjmrrcmya45wOaR7O
qxH3HhbKfqgvrWek7CTDDYaQFVkm0PvMjxmWpIX/ADBMvTpT6PXMUw1xJ7+Pui+8S8QFpUZuFJgp
iAvPtN8JI8nXRGrPRRKEYZD4sF68Bb2qkXEP17B53WeK5yra/zl330FHkyLjfiB6RtTMcnyROgzv
PJ7co6EnN7KrvGMyFuJFsJXs2VppSMICNYufo/aOOJ4n/vxwsIkP8sqEOjqzquuEz0SvzesCqsdD
44etbN9Vdwll9NPWPNhWs49eOsxb/UJnWxvd2Tuyq0Iv0vAPKkAuBpm/NqCr9YYHiGtEr4XOMMls
QPRxRy1suvr040tQtoue4fI/TmGlP8Rpth01tY0TKC3ivnsJipxPFHE0JmIryBwYN81Gho2+GBY1
oROZ0gIKuuBPtFBkkdhemZ33eMEJi7HDny7UNAL8Tjd81sHrJHp0VDaHZOLvn/qk6Yy7V6S21ZpD
aHqBZeutZaOHZz52TxepO5ilqHb+sVXh+P1naOWuS4124VZH5Wcsj2rM7oW6myTslP/qoV80kZ03
M8faFzKIlCtK0raploU920/a/hrQx5FpA92Z77Kv/ByyeAkwCJI1ezYESFXkfg76DXaVbummbOlS
Itc7ebWa8WvTrK3KJQk5OOnbMnAVFtCj3AZxEdoaKCkfmOixCALAz4nJilXZA3eUwq+aDhhAL5Xf
y2pkQ+zq/U/Kov3h+iGK8hJtZ9l9p07JEUTy5HjLIDJMDU2IR+1PQCeIWpPhXnvUtCnCWEtYJFk6
9KAnBezbOsoacxLeMMsXWnoxwpXy8utnW1p36sbjAYzEnzRlCozdkjv76dQ9EL7sqAPPZffZ8v+d
MJy4F9vhCmpkVVzNBrrkWHO3L+inzFRDk182O6bDXLwT3m8g6nvk6iwmtC1N0KodAS3ZOi/RhUVU
JGo5V8KPKXiNEpI9UBSAdb4atTpL0/vuS+ddGLIararKbbUqdaOb7/OszhEEZBdgpROihyl+0+PV
94jtR6CsNboJHQs9UH18mUDS6fy6cUWpHBeL/RJtNVu5Ha5gDFUcsgrVmNizDbJhOud4ApjOxSLJ
MUegVGy9Clc9KW214PilHL/VXlvtMqDzHmGgAx8PFd6yH3UjUcW/GnCrIlnms6dU0liZPgnAMSUy
Fd5gjE5wzopgh97POAKk+tB1Ej1qqhjMzmMpDSm+RgIjfuOzZcNSGe14bsYRK91nHz2SPqe/pr3M
tftj+enwmeMKmBPfaWqUcJvUl33R1nJr6ziNSQJ9XswYCj/et6kWKHNI0FbsVm+8FDNAqBrR4Eyc
DGK9GCbUIU+Ls+/5mEH63pxJSstU/gdt29M1FTIvbxh6A3fL/PM3IiS+AXyLQpF67/B5y+5G9GEQ
Prt+NP4Vj3pOff4X8URJWxq64YmQdMIp0FGSj66yqjFz0C4fkhKoJhOdLI1edMnfPhovRVbCP8Xz
UpYzT8SZyD7Fgk85gQ5f/Deq+SVcVmqhcYIgLQzz7B9KZ/uUiOq+KbpTEJvSBbSMCFRWMpDraSZT
QUOvUGJGNC31duPqYBdmp6QOPqDzyj1WcOJsqoc7V0zIa4nxK2sR1HKD2gaBlv0QR6k+lDlht4sB
eLvXHnz3gaRIJ2LJab2T0JeJH09g0AE2t3SjxkSdQUydXm2r5vIgrTBKFwcz2JaqRJM2lYTPl+YN
QjVjCT+L50WSvDYCRsa531zx2gmTHEWFf60HEi5Tm3SlLVIyXUcA7EdYN4IwhTbDz3iW9N39pO5i
8cygtx7lJRw2gTVenvtU/CU079AA5os3mHH6+BOwPQz33ny+HQExYoxBLqh1qfXRJmNa0Vx3BVmi
WwmdueYOYpj43f4hzJGjmARN/O69jxitnbiRW0VJKlJDcUfK40FS8Qtx1CWjeBKzSdHDpYkLAv/k
NpaLylJOzFE9phzBc3U5LaA50IQ1suxIT3lsse1kdYXIc/c6KAjTOtjXGcK2prPhSQ9PsM/87Cpe
1fOEcOBp0fRtsjyjNkgDomMBArLbLAXLFFcm9KmgxHEUi0iO5eIQ+zRFHfcA9vJRLWlJd9mTSbCg
BZLW8X+Mo+lB6iJ2Th12fqLzroRVke5xSLE/d3t2+YoFzA3YhYz9OoMvoUg+ah8fUHs5txHmnRlM
JjrWockLIqlqoLcdiGmUUT3SfbMbWMNnGkWUxlG5nNxVoJyfo3KBKwgJNGeOCNJvRdS4+PXRk17I
p7H4l75PfG4zdY4BrswNUat4Id3zGEgeRpkCWJPfLO9mbb6oBPoYTzz6pSR8mEde21Yt480hmZIN
oi4kBLKuOZ1/L20hz15WF47VbjNqWK1xJGBaUsw3Vt7BuKsS0aZKOYe0n6wJ62X1+m4qh8m20c9f
SUCHMhn2K0Km4k34ia/ZdKDnH4DI/WtVLKFlHfHf55Gcjgs89KpDaLZKQ7/6rJgTZCBlD9biiZBD
05vOZrh1eAkV09u1GwfaC24+qHHrT6YSO/OY7e01WHTE38ebA28o3psPTr+CnDFWMCYUo0XPVHtc
zlL5XDE8/FXjAfG7VYZyaxYSjpaCPbK4G3MqMuNTppUXqM+amlGz5TqJIDJWGZ96LPwwBfFTzrug
JsDN86vvILePnDDyoqlNj1Ewgm2cHxOg3Lo6zPzq63wTzjnWxudYWkhhCIXyCIgv23TvQNVthSWh
zUe8eV1RcyhzJI7V8degI8AIzPfxL+uIY7sJHAdmisPaH9Lovc6LGFtJstJjEikIXQjslTxVZxcG
6FRkSs/ctPyQzJ7iFW8Zms462UBZCbK40E2SjtcuG8bVKUkzh/0DS5v0poiL1qiGSZHm9BvdvJnB
Z9NGVEDxWmEzk9XyzKLUFvX3Px/+k/On3mkmr36mpGGa+ERCx2wHHR1rwfeLDSN2nuT69T8MTirW
nta2e/E3PDWnJsyqlGQR+7OD4/Wkcj9JlPAD+0UrRGmE5BvmJUYpZ9lZyHOMy7DdyZ2LHt8Hw56n
o95YLFKb0xQFqSjOJ6ScrPtNM3zouj227IEbte8/FEdxVLkWBlBAAGJMgVWTQ/4F4Nz5HsPNoU9x
Ecwiah/NuPHCO7A22lUtmd+pCxZqANjukgVPzJuukb0itA+FM9uoO4tnpzfFXt5IC7YuJYEeN+u2
9C2XzdRgy/1aTcCSVirolCDufO/nbPNcR+EUSaCa2uSJa5d5/yUuSoqt31Py89ftTSnMyQrUMYJZ
f3AgPluErm/usFHkCNEeGmzcn0BUfijn548NmyByqJZuYwgzqqDS+jszv8ltrKACk5ir5PIDuWtf
ns99JT/j9yFLKqLSRyQcVcUDPRM2hU/jnj2meMmk+PGStOpW/RLyeTGFt9sdpcgbRJIdYdS+R7Dj
N/yemHG3q1okAu2IcKjGMlH9aIln8+MhfL8GpjfJWBNDp/YvzFr+4okBsEFDzy9nofhsSzzppD/v
r48xDCSEV6yoEihvMMENzscxinD6t8rmYcMjSfGMZD6imiXepfSWvSRVNwNAZLblvBGrxJpkTLOj
q+cGBhjJTP93l/Fg8rYTokVylzD8yOdO5iEkyoN0eO5+OnfmLpBvCV8+Pn5h+Sxfqh4QnmcrS18h
HsCuLzguVKozlCxNimZkYruYneA+c4FjKdH4i7NbUei8pvaIJ+Yl5ovMRpLVTLURMveL5L7PsX7k
BTtwsmuB3VQoYe/labrecqeklsKPWJmQJYx9+yiSbuEvl7+ydjO6k9Htj3poOfIkn7p5OCnXnDb8
BgLX+EEHhlh2eM5jr/D8mZ2LYG4LKturCf5hhZDBVyc4ahIyXCNH6gtGR8/pEIF87g607Ay5cXop
qzGVR3mywIUem0YR6Ug31g09S0/kgagm/d1qBG8Ph67O63tTk/bnk2vYtBb4pAl69Z0IYvoVAmNX
gNXLGZbqkGVOAmTQ9uHRaYZQstFiXhldUyj1ccnd+39YsxjjxdSca7YqHfZvsbL53/JsWHgHfeAt
J+Qq6Reqv7Of5wqsMBwnGMq1hBIp7e0ob8+tGd88w8C5iyd3pPjmdqODP9zLHg5/kYnJOADscHBX
uwCE0Zuz0x/TxV3otW6HK1gF+H1z7R4W/w808Mj37S19plG77mAnMhP+gvwwjrDzNRpBnfS5ZmC6
B0E7eV2P9Ik771IUdU/b0UoFw9Ui9eBb1Q93ed5Rj/KZd8ciK9tDr0ZtxE7I/jCsZsctJbJaduBw
iXFElp+MyAgaM7i64aI1sFKEBBWs0oS8zYPIvFHkWnaqmdjZjnj8bbEy5tPZuvqV/SZDyt1LUz1b
0/KflhttXyUFEkXUjeSEiXH42zh872trnXeWul5yj3pjXol/ZlwC0frzYjQP4BS9kDJIaKC2BKDk
JI1n8F/6a+SmFVR6ssBJmmNzw2gGr92iaW1nzVPdpjMh+S6rwPhzNaTlvRj7q1ZyMOvY+O3RAamp
U1kHMeuUZNZxC+mymWqaJe9f7ecb4JwktXPKJyCoJer1qKFlWaA/D0ksnYVeg9+nYXFrQtiWlymg
5Tepg7zoYnvwDrN6KzmrASw/im8MQzpZtBrBPF7nwUlcb62yzB3ml29VYFb7W03WiiWHHfeQE++r
COC4Pt0896nvmw8YY07uOZE8rWYAiAnh1tTuUas5v08RwXqxNsIeN73SfXzr+9hIRlFisslUi3O9
YhVI3XGLcKmoQuobkdYgNVVufi6T/7aKs5nGTy3CiHuMSOiBGatx7ykB7gwhRA7sD7EcX9xyVooi
yCf8UwTtIdoy7ICW3Kb6E6z3j05OuS1bGOyEIJt7CzwV3kbc6PSUK0JCtwCnYdR4zj3C4kibemNH
C/wx9D14J0DN0yY0MG7orFWO9yM3nxMlQHGl5OQHQ/a2WD4NVdr5LZwo3R9Fuv9frKoCUR7Hat1C
9p5Wyh0TUWuch6QsNBQHnouI83aP4mcXYzdbJG20JveMeatqgctxDMf+i5/ZhVIxT88G/nMLS1Im
3eliTbYhZ3wTYIFtbQ3T3TKzldQJiy3Hv3wSxsdug0+4I5Ksv90QzzGGMSp5SBUcz6NQfeH2UE+m
azaq23amYthA0SAD5E5xgi1RczV1WZtvRuFzhRcHtNy971jp+KwcEvp2WzaO3dtzJSujqzQxZ865
wyHcbCQfoPLLRWqjGi7T5B8lTGo+9nwh/CHzUVU4nJLCF/PFAOmReBa6lBR8/+3Avx1z/reWlI/X
KIPZeGP1lkMtPghxa+gnyPPSpI+dp5/J+FW6+JYk0bF5yPc44xRUfp3hlt5xQCF1Ehu3mTy1JemL
hmaqQogKCVa2+/hnT5e9tU536h+GH8GP1cIvTAXCBzrKfUhg+Qx6K9lOEp8pG6ByikjZYVP0jYUt
7hvl8RBAz1Ns/3iRpejcJ1DDjT3AcdNfjD3CR/E8YI+mXhq3dWTPWDCwQgcSgkc78916BaHUX4zj
M6WJFuGOwo9ikJL8IRT8Yxqn2y72wPm3HBvsRxNMS07VJIRkYDFqHs78WcZQz3I094ktNLbhHOet
nOpkqA16IXlCSm0YtLbkqaiz2K7LYIA89vzEM1/Dkhgum8P5ls1x1KLSV07t7MAJ8OyPWH3/rR9V
IvpecaUS+eK+4R5OS/3mFsVzQXPqD380ytpMgmk8pQEgY8+EBIYGmQNsWiqk86q6Uf3cji7WF8Mw
BdSB3q/0ckDVtg9vKGR32pxvZqO21iqtNHA/lz+4WeV7Cck3XyovxRUdqkzucuRB+Wcmi8E+WsEk
haVGCQ2rPqEdMFxOXIgdLiNOUF1eM6QoWD45RpWnj1p2qCWsKl8xCMFoMZ65388NSk3p7cb7ircs
j8Xinc271OJ49nJVxoQa15bnDWmKa3fe0QTFlBfWLodAgCg+RbPxTvXboJfymYJ11MsFnqa+khiv
aJZEoiq9riN5VvfTPrWgxV4Pt1ynwmZZyxeY9Zs/aI3AZ1HGCcQMon8vS/Kmero1o4CCaU+/WZsK
ZP8XGZS57KSe78R02wGUpOJxtfnoDKGTD33v6DiQmBh5aHu/gZl4hjEzxignawG9oBUSP9V/ECdF
wkSCVINrYu9oSurD4jvvBRP39xfLbhOrOUiWvN49YNzn3vSY+Y1ujpSCKc+WCtqGIFBPtjpfUBgQ
nnH3Sr4oSsuLIbgI0Kqax85mNhdwM9Kk2vB7PCsM6I2Y4i+ab+vYYlsBC5zWvqdfyUhaE10Uja5G
l5y14EVVcclmn/o7As9qYfovo6Tdtl+/F1vBKLCtjSmbbG8IaqaRtXgRo0J6tHLqyflgQla90uf8
bz82IOzFdfphS/s+J9fSiiIf4JhyXNMnyfJ25s3QecijDIzuLlCjK4tpQoqWTCErechfMrPV8qTx
2sENdv0b7DDKBMwff701cDNvnaQVSanpo0NYQt6Bxkd7wmeNbAwNU3LgU0HN5jsPCd0hRona4KbT
APLckHT4eJc4V+peL3DY+biJQ5rTX4CkaV65yUEHDY32SMEc94M+p3+oRrJkmZzDYY7Y8rZj8kG5
pfvcft8J5ekdZbhNTthMrenxnZ+l/8veifRo0BPLyrV4j71tbpbUGhDwK4vN7+4NqHX3CP1uPl5C
vysDerPeJp0nJOjeEpthLx08l9zkmZYiSd8kUmAF4omTuq21VZlm0EECva0nFrj1tLvzmZTCbtpw
yqjh/6YLKLc/N7ptUKz+3KTnX04Au8PT460g/alJaKMEKx+VfhJfzD7lqtHt3JVHgjywnpcCE237
iOSUWxDfGbyyg3gDXMqvERweQ8wN+nuDSyLI+wfqq34JZAdMl00+/q5BR+/ZaqITDBvvPD/WaoBV
x75bChiGaBe/CavvuIEMYW6CaKnvxuKXPQnvgtBNNehdwDeaumdeC+Fnqc9ZQD96+EXzRukRw8qA
YYCVlPEdy6KZ0wtfHjNBGxIGICXhp3SnKttSj91L+Qn90Uqzd/eKWTVzN8mTFeWkmidFBx7owVrj
Wk0UbwCwfCGhtvbqsh42yvBJLGglaLTDjm7iTljHiGRUm60/RvzpmLcvu1vaRVGD4SEoQD/bV6Yx
wIGOZvilrw4yQxVtUI4PD0e5B6HJmBhKeOZIs0iRUM7pljeSHoBBbMzMoXesphtdMbRPaCJLxc7h
fBOdYROLAx14wXs2vWG2ac/fi/HmI2F3kogsYza9Af2Whh/2yBppZcRh8ubuAp7YPf/WCx8RCgxu
McUeBHPYEI1OVjIx6Qy4bpdBzP2DEUlLd1SOOzJk9szowbxc8Rtxgglle+/jkvZgqg6xIB7dozeG
GL+ZcEaAke/aJM1rECk9kRI0fe7b6Ij4DMYvJRxlSWt773PryuMmbA4uvn2U1Vl79eL1kCscwyOP
syxwnHgcbIkEZGJ6shxP2iEC09jnz71gbp0uG4Wh97Z5EuVHYj/I37jcaEvT7GWNQFyFt+n/fv0j
SJ+KheiNyOyFfmi+88nC2GxUPEghGxOOmKbJhZA5evydvHEMpQnYw9HxbiqGb83KIis6P1ba6EXk
WnNatI1uOdJxa7M4S185DF4QUIl7ky8W6K8Et2sZ8rXBmDTXcRqObccPSpABt/WLjE0yqR1StcSY
yiM9EDFV6Gow5SLjuVf0wZVJuCpSNaEDu5g7Ol/sJi0BNvCsPIh4mvKIZJhcIAqM58TLSqgsnZXp
UGbMBxFMP7I4gyuJQNmxNeRhpgttJ2kySKfg3MuB6N763Q/wq4wCTCmxEzq/+BcVy31qykqNWg5t
vMg4MPUlIGrE5CDbpSU8PMvIFKQMbikH1DR/vio2Jt7McSdQF+B/AoLkMWQQyI+AZD0xzxQQ5XlA
UVijmxiLB2QYyJImtTsYdbfYvKorhCDYGL7GJNd1xPmJk8tZU+Xkb77+JUY/5FpLrrZDLAKj+yGi
EP29l4ByrAT1E8PYrSAu4cz1EWCDc55HJv8scRx3wc/gzcPenjVf2DvbhhQyvSmrxa+b3eD5HeR5
hFd338R5qRIH0FvYkLEBBee5GCv/ex16wIQllx/LhnjyolROiEPidmLDXW77UjCXKMXERoRo8Ne1
00hkBdppEoWqcLBJdp4yv+/Od3NKqz2E7KJtXMz/+4SnFpr4wIGQclrS8p85bF4wNVn0gBYR1I3a
t8hscSFtINhzKpxcfjV4JiMZi4/aObfxSXyyLD/X8vVh1XF/60GIgfu0Xec7v4v8QXd1NRypC3xa
f/fx3O2jDbCB5C+Af7aZbySNDupnQo66hUn2SxmA00nmXuStUzzBsjXPdKfh4aY/i0qkY2Q6SJBJ
d6/iq/E5PMCPUmGnoqLstjVPNQw1nPLzuHBRVGeOPLvQrOQfuC8Pz6adzo9lVc9ofWN3D5pvsYzy
F9kNCGpatlqj0/QNghSqRCEMlfq0N/7sKOMF6gbhH3x30zLqMy6fP9YgQy4REZWOXByq5syLUpkY
2WkfRT/HpbLm59ic/uA51Z7WRj847eDxJRO5SZRwuoBpI8Ts/qyf0iAYfwS/1J4xmmJZVDvpcToB
dhSdw11yEZu5zdFwjMQQkNrY7CPv/tzJT0z0iC1x8QFmGpv2+lR4mRXyXVmyBYBO0gdFvVFXA3TD
L2GSSd5s9x+fB+MT3agX2kfj3K1gghZaPBgaDNVVs+QP9J/zpqwYa3Idm26Ge5a6bpGDvN+4f1vE
dkx5vdw2kP6R5q4tqyclnHfJbSUHsTV40284sRsZoWg4wl66Ov0Ke3l6dB4POTop6j9dBBcr6IBB
AZMtuaMF7myTyHRy3KptT10IxoNKSPoRfqILfk/YKX46SqEIZR9jntbBD/bFLeWXuxk3C/Kmhozv
0eU1Ot268q0EcEllvrlyZYhOpwqlsor8FAi17Bdc+qHMpKbGVnAYzIjL0XsbS/DPex2xtGbhroaU
Njg33JBHwibkZIvCtaduRuFsYshRAxq0WUIMo47SohYzbullTqbdg/SrBPBmy2BA7uWQKQDMJwYf
Fr5/tIU1OIgfZ2mhEUnzZUfEncsJDCo5GHMpFa907QzhSOx8qA1NO+jBWE3HDX1nQeEEqdMvyjuA
m9vTitvQw2yocm9Z6WUvolxatn6mdgauMbivo1ZE5T9LKvEQVxxI/1QLzQroVdsXHjZsUy6MPUEP
O6oXIqemw8isaMdVcRNEfC4RyU9rBf0+WeqKfPYT4pal2Rh5XKWZ0vguKny0ks6bpNIRf0mmmGmX
Mz28oC3JwSIp0p30dMH9qs1kqRqcYUWObzG2HrxLaZTVlBkblMky7XqssbF0X/QacYnPG9aSm7nG
lp0NxWP5b4vXfe+R3yTX94gDlrgzDVMYOdRWnLyDZsyoh6qm5SOMxHbnuY4v0zKG4KZ/+nB7TKu9
flHmCoZlN5eLCIRFBsN8FFIXwwVhls9Iq55xkG+2MTXKKilN05SbviYl9V4L3kujCXOCmLZD04b2
Fy/iwIKFz6RsxH3q1LvzHIRmUsysnxtJDHArujN3R4w2up3T0h0aEGrI0Zcmubx/8dYvJqxAJ5ls
GVtD+8rtm8/vZsIyhWhW1sguOny8Dsa0rsYufdRfVRjvHMQJD4T8YKdA4wPGaX9LAGx4ZcCIHhdw
bq0/hakQyZUoOg9+OTtJberaP03kojdYXfrI1EX038sbDhxlTaiEVQppN+AkK0UQEj1U8LpYg90/
fDpz/m/9h+mAqHrceQcs9YvGsIhSWwKKj8Wks8slU/uMSfKDom6rLnNfwkm+c3UVT6xFeEFbTklU
MemVxD5mlw+IEQPFmGeICLiQ+RUPpBHAy2+OvOPt37GwQJQ3P0RUdpKkvqNrB3cDH+l8pfx0qEWI
IrJwjf/1lKjyq/HD+led83iOY0LQSW4u7l0NkdWMDc4PjqlVXD3rwzvyC1i8ZiQL9RMBjqWbiste
4qRWsLGEAtUN4telFjT+eYWa3AbSTuw6Wlj7w85xUqxIZq453nY40P4WfwElQllGw612a/TXuyNi
wdaPFak3H+Imm83P0+d9boOiBQKpcihu2L3gwURBpS3HYMk+pxIicWKVz/TmZgfNq/ILVeT2Vo4E
epRmoSTXcVHFSCUHXBNlricoHzOpKnYLP9V34k6whl64EVaV981Nw2F6iJdzo6Zm4SOTFgcSJ/8E
kdN+qCCm8Zc7u5WKhtnXiA2GwIEEOqWoVUGudZVtfQKpF/O6iR6FX+tJCtTeCyiKsFSiHrU8cmJO
SL+T6mKssq94pESWUtPEApXQrtKlM9CcEI6X2lbkhgHausZ/MuYHOSKWYLn9hoUXWIqw9LIxb5Pt
5U8CbxyNdExmAZF0sDkl/F2cecztAGq4IaVUJUOx7bHJF6H/Au+//mxeudh/LZI5zMMMgDw4dEMt
LqSkbeMTJiTsVqSAvwohtfszBtvCkWL3/k41Jm2u6iclOoOfqlxdWXKohFUgjImrGFyWbijLzCst
aNb34H7ZcW3nHuMWL5QdsIEVHeoM64g0JwCtVVDdhGUChU8gNUOaDFK9igTJAgvLOOFNT+hOS8Wc
DGxbRlggqLzBP+GT51GonU9SCVr5EbeU+ZNsGKB3acLvEm+gNoKDxxBeDCejxoF8tycueynaaY76
elsryLAkpgKF/WXnuINECPZr8Rc6At0cygS0p8M5y+RBIdBtj7iyI4R5ba3BYyelSZhw57DJOWzy
jzxYIM5z7kWhYdtHAEJ1td4s/v472I2XupqFreVEH4dh2A88HI9KkwKdUKyfPkWffVvvIciX1TDQ
+I4uxnWMBabCV5UgIBHSv9vjQ375HQbjw5/85VdImJ5sbnIPX+RhEbK+gec8eIyv5zkRC2ZjczrD
tCQ0bZqJ/qNKqR3W40Pqb7h3irjk/1wj3IZm+Y5j7wDdt3zx3C1CLBpi5BXksudYF+wtN7X1NBDI
j05HdMorvNtpnghkMVuT7MXLCU1Xqh+2LKMdO4Ov39ZGzvHk85sLQblH8+icjDGTVH9a3/31t6AJ
QP21MKVIJlxYGNeKUG/Xft1KVHLDG6Q3moBC3oddktTQg8Pnv4PuReBft1pyvowGlb4fJzsufKUh
QhbBMTOkxeA4XRSq84ZKrA4AEBm/EbrLGwGxMklXRjU9vd2NEf+lmgscgz4TA6pqF8ZfCDFp+x3M
b38gwLI3tI42uyPx0ezE9aV4mjyLssvyrZ44Z5xb2mx//QcmqCGRdqK3wG0repZeKcI3b/jB320m
gsPv8NrkOHhIBNXO0KZRqEHwE8MrLmigDsb5H3cscM4OvQHbZega4kFPjgK4LXUCTVxQxvJl2NxK
I6HEBexJ4rRtHrVK+KyCfQB4fEDQgSL54M2PX4RndRK0JuZdSICYGu7OPkBD52RpWrETjs2L6Xb8
KdWEaLO07QolKTRXIIk5/fF4wXw8RhkefXmm1BEmZuzKoa2H6EYlTjepuN4dCyan08WMmJHTfOsO
Q+tqF7Ln1l0LFvpmwPBIcQIDm5yPk5DXVX3mxs8ddaztzrGiiX5IPbL9yOPqvof9kYZ9ciwblxhc
4GCQVjLz1SWory8J/Og53ynaFB0/TkUHCYWleIHOw+elQw8pk6SZ/szzUurhcBGG3dcVurUKyde4
CLYqFvAuBN1SCQtDAq+2KrsdXje6AV8Mh40BQr7vPgtjuB5E+GuP78GhXoyMe0U7BZQR3IGDWPHU
/0aPw4mUN8CMPizgrmHefg/PRaE5nNhUufEmy3WufcR6USXue7O+xd9WdvkAOzyvNMAOG9lk2kSg
ZmjGC3bw6q7KuD5w5jko+XCuSF7pWk/SmmfsT6+s/H9dUlLKfZ6NNOa0oqKx1rjZc9/e6tSmOhRv
WkJJJAtEq8CAOueE6EStu+EwMLD+tjQrv/QL4z0m7cupV6w3osjYNM+JpEBvzmvX/d5JBW6ygpL4
kgIsCwb5FioQUylUGeFue3jQMMAJxJ1tx6CVtRhvM22yMgpbGYXBr2JARieX44HvHr7aqu2FKPAq
1hrdq3SdCI3dpwAP5rDaH3vk6LooZIeQnVsafsUhasz4kbM4Co1fRiOG4rBlVXoiLTDmLi9KqQSu
R9PKLdup7X8Vlo6b3RCT7keQ3LYp+DJ2Fp6ZqSqb6API4YWZ52OYWel5ZqREee5PMT1RwaGQNw09
d8/vGap+DaSCYCk7iThLPy4VdUcRtdbDR7gzNnzDU+uXBShxy5xlNvDI4SWXOpqhQ7Hq91xGm4oV
grDxJFRvjdePB5qreVWW2SjblkFawRGJuBAC5G0GLy6wQIZWskcXEHIrUgEYCpwx2fHseKRXLty9
C3rAeCPc/p3wW+xLluhCtkmPANuPQUK/SunKykYeRv/Vd3u/F6WBtIlsaAxsEQxCOdtlwZnfMW2g
/w4z6gXJcFuVOTnqJNGORchu9SuP2dgVsXcAq7ROmqtUYO+/B5Os2B8hm5D0L4X9DtOy9gdzjjog
oohQPITHdqzrKDO99aDrGltDs62x+omXD/F+4Zgns9r/t2QRBg2slf0BCUoErOONDU7wz8qoVAYI
aLrskGK6pWKn+0Xxy0xH8HxvVgpsjC2x9wtdDFUVP8lVIUBcdaNge+Aq/XJUCQZ6mVLalrD3Vl9y
Bgj9AzGjIDK3QjPUmFcMYtaAcqzEeiCMoFF4zk404Zd7AXHe5o1EmOmv6sn7umX1zYNpOJiI3yWk
mlwu/R0ZehIQLw/agx6vZSG//DkXC17YHF4zumDPpTmYTQkgKJvrqArk+osC6e6l5p1Qbta3rJHR
e/S892v2aoR+TXHH/8tXmOSzsMP+R/FRu3Gna9s2DOIvY1D/lrG058lFKxKTbEjqKoczEfNtIBIL
fFR9a1e8+TtbwwUgo7WMxCXm0nlgVxg923i86A4BXLCFcoWy6M0gkONn5wadL0ouG0HFZg/VDAlp
TEtejS6b8H+icS1V30695KUisx8TewUwCiguoCg6HHcaze8Uaf1fUyXiA6JezK4uqKfuvlY/z2Oq
CIJL+fRf+TIqLqwhLwYIv/rmrkPvR8+2Ptc8WQn26rXQBtvLxj+SR/LtTlu74rR74CgsUJx4UHRU
O6pozjtid8GaoDtzIXk+qNmb8c2p0ZO/YOAqqM1BzCay+LCg1kK3TRng5rrZOOJKTDfiGGD/bxvm
uZRAN5ttM8yq7lXDzs/eaW/TSIPWZkZrFd38D8J8pJ6bLkWG7YENRPgcvdSyMevzmsMZOnpoILO6
ShQAy0vbVD99W147k/5OMWLvlpihs9qOhV9m3IfFG7Q9cMpZpz17hL4eedaUKb9Ef278KshWVjnd
yrauP862dh3HaiS/b6oFH0zGWCDSpAs5iabXf3FQ+RwiTjAkIDJh/t2WmZMHxlW9tdNJvALBujwJ
nln5HIKqQSiMkbwaIl0oEdbv+cbLAmpT2CUEPwd07gYfRHd6AOeKkipdkQ2Mix+vNYsecAHjxgn9
DtLnJNYdz9T9UjTBSv/WTmtU/nrr0qD979UbHb2nDW+aYaAwvZvx2ZyfKlqZAtBgig27dwqg72X8
GeWQi5ihcx1hXdY53fbF1UlsZDdPzKsH0mwxlqyGme1JUfMCJEqn6EOng6WpANOBUACeW1E/G2Sf
lbZpJlMqEmNjGlkuPRk+HfIkZx8wqLYWWJ0+7uked+BH9H2JlnV3erJSf26J15GnAWd3Oh7gMmNL
1U8slvF0pT1jW13vAWcpfevur87ea65SsW3X28Nph+TyXDHpR3VrF5SNuNUO5m6WSmM+7+gqLCeV
/BNg+YzXNfOTWRCnXbym8uuW1o0NL+/R8yBlOF77k3Ltpe1IjR/BW0Q2tEWO2B6hkQckiK/zQzHO
wu/NHn0bGliXUorSmSDemV5Ao4XZDv1rgA+I/HxRCD8fGOzyfReq9cbmmHGTXp4pBAzpw45OrX88
TsGt0mF6/fezpotF7qacoK4L5zOMq3GPDYxsotIUgvdown+F5+DuTN8cfjVNo0tvtnUvhKE5PtAS
H2LN0/N6Fjcy2H/NHbw42sbWK2ixqAhqF3ZwO6lArMrNRNiybiyNNqUdqoI6ZxkZnT+IfCI9tpEU
RJ48qpj/tsVBIC68uzAWIaWawn8p0XrngBFI2gVmDZEM2NOCCUqsR+D5+C9tbDsUoLLRd0leWbJu
vBdZuSRxoWd0wUJSEV1lmgM62SpNeKZy4WDCgs5MXxARdbx3AkYGa9WHTbH77ibr0pr5pP2wk2Me
4fiZMHs/D7n4h7Q6Rr1F5TP6h6jmlFyfdAb/8nqlgFixeSzt2EHjbAkijOxqZSYmF4fe4WyYrIrH
qj/rMAzY958mnOD+oP+Up3BmHRv9zPPcWtQpvyujTeb5tQ/yLu3XkchNduRNVhXE3UswyNvFIdVh
8d4BhFrd32FNV0vPFtRvO2zk3HR1iTBJv9DvjOXt1St4tOjVrgZW8StiU1qBgvQfZik5kHtVJLeK
d6NWEwLstpJDpCrWrkn+lgpNEfzdWCxmr1ZE9z2kkUSR3KcTsMyb0IHPGH9zfug5JuJdopYzc81S
SHoZbQPgrnOeSjuCJn4TIBHXM4/NzWcZ8szR0mh8flIbn9Ozr9gKzhrv1qNv1TusgdFeXNZ278E0
IctDGmXdlVSXKWktYSZibslcmhdp7Tr6OLLeYN3DLU5a6ggro4pDHBpsIK1hhNSQKqXEHNRwrJDq
OGDXrL2iCrLakCeMJMWtGD4XLm5UawkrrnZIMNBkumpvETMELme4M7Kn0uhoOu4vX4HDGtbDeUjc
PXriZb4w+dD9YwkxXQMBQ55OgWcwnfE9lp8O4pnZ3009hhdBORqvpmERKNnsQ1wumeICR5MnQ0u5
e5rUxX7EO2TelxUgwlTBSkE3e3Gknz47Wda7Dv8Z2Lallm0CpIwb0sFUq3hmFfL6OBp1fO7XxNl0
S9lhzeSrPYI+R+t/YyqRIMPqYNh+wifRhIfjsPQo8CPdWTJusPn2z2BLjzFdTUDhl1SBz1WcimVV
HYIdacmu+fbyuGBJ8pM7xgqbaNpM5/dVJ/g4xgnZZvZxTx+QDRPhW0bKap0/51bmwr1V08B2aGJ8
HNnV2uO2TTX2Hxx3gKW4iJArIVnawTi6sWtFLOIqIGcOcPH/Jvy6wuVPgEcugn41yVWsHh0zgcvZ
btHuR0nKUkEfiss5/1BHr3cLs80UnfX4cEHx5/8RiPYAlJzd8zStS8XxMhrEy3gJaXUviwRQkjCs
d1/oC95Lod53AeeVZteW+f/ImappewWJvg+n7eFA2SbcFLlWi9HsSYL+vcyUVCevI5hhbxD8fQSS
PXPrC/QCNA4SzAm8FMwFkH5LfPaV6tRqpZlS+UrAT0NuS2bWayg+9CnurhpDLPYK8I7cS75Cjtmy
QA4X9wXrUsDtXAWVGZaSEBZxKdjsYdpr6cmqvg9Dq8S282639Dox3fng0Rs+++26aefo/col/Kd+
j5q53LPOs+VIPSC6EnFeQHQgjeL4OKuO78vwNgKmlzvrpSwNRSvEqMLdNw+rd7EqoSmKhURJi9b5
dAybjrBO+2Jv6DClEvFRZIpbYjK8eLLT/xhBhS7vZFp2kj/eyOby7XAgLqmLYgLgsBcrCBo2ot2/
gDZuBHaGK00MAKZLumWy8HuAEYbxndzfXjaqiwvmA6oWjFSbBmhKVNRuiCGkhbYDz7sQAmFuEnx5
jZ3AlmBoVLCxKxWlzIrlbNmR4dNMjPxvz5ylZroRqAypnt7UY09ikAORe0o34B7umsHlMc7vQNYx
g2tZL5D4RnGJThZBjP7PzJGMl1ddh+hOoXqp2PdDyxqzvwRDdkEX/uBPTRQInIX0khURcWgroWOd
apZuOctv4yOvid3fc5ODv/BX5OjrQCgl+ziM4OrbuuOg50G/58LtDZChTcAoceE551B5hc2AQW0d
4SqVzMZmUUExbH6L7PVpAcu7khdkx86IhArj4u71B/EV7nJT8gRitN+1ISDpS/MZF5COs04seq7c
it2THO+wFWVOq/3Dvsk36FBq/w49W8deLzjAEw/uecHgYaeI14JDFrmsZwtyySAaP5NATxkHKjKy
eWEt6zzRHbkeo1byWFe511+ZI5oS1t5giBkNflsLuyBl0k10cXF1F/BXms/xqMFcoOP5d94L5DR4
gO+5DPoaxRAYp9MtE4muCZdMy6djTwoAkjqu9zSVbP648QySWTwF232HjaqkgAvhRBvhE5Gq5Geg
T6aWOShTFx3+hbElh2tT3/ki+ON2BF0TC32nrXKuTN+hkm03F/BfW4amzgLH2gfJzsxUTe0qdUBT
Orl15jx6TTVlEdFKSwZFaiqTUr0hXSuBfBj8cvYqzmD1n34pZUW4bds87EPQ2+8IDbVPPVUxP4kz
gRa4BMJgYkn4NRL9AB7AB6xSKEJ93EpLqSg/9ZXb4H5W/f01ObdQTDqPKP/JB0zpPMvgEuZK2Q8Z
/pSHkCj6RKiXb+bjQSP4P7uxeY7l4KGpYahRyBaVPRFExW647ZopDhiRSPtNow030Q02j1heQqrp
GMYj0FPwr9Z0j4RHGBHo1NgkJIWy98S3D4wyyxNqi+T2sDRWCapRskPosEwxk3owBehN1z/gv/jz
lKymoB3btUWrS23ks+8adkKALThGT1irucJkb96jSWFv5nChJUNMHVF7qMtKBIMr6hBUxLpTKJKL
sfBPwpcPMWNev/OT6QisEtl/rPKgGzfrQZeEbga0Ou/0JxD6w/2jAzJiMHHV3Wp0sg7MTTMLQ3qV
O4N9jP+1x3QS74vhNt1MYNAlGtTZTj99WN6zFQ2XKVvgwiEDSYhSstjAYNz9Rjix8UWmBT/Iqp+9
+u1m8DrAWM8XtNGu/eY8t0zoC9p6E3PtftGViNK0giMTRAseeFj+E0AHPldmX4saLWIgEMzXHtoM
oO+mSwQY89BhdS1CS3DxztTj5HrgYF/vysxIUZG6QHWWQBGfieUPXXjGN9ttAwRF7nEl4mgVLVBz
SRPHtxC6RVWk+GuciQaSC5L7DpPz90gtg27N5xd0qBN9JGx7Amvp/d9CJcr7ArM6ODP6hpQTOI/q
P0NMm1bkXnFfh7K85t/ztsjwhIid0EL1COPk2CjUG6sl5luA7qfHQ9RM60EStSFggSwyKAyOqHsW
x+4+X91vYIGMj/FyHhnmXNnU60T5y+D3ag4ZKTkxeJfm50FBIeQQzjxrLZmkasuwsbLLY3KQ7Kxw
VBHjgS+/khzRB2gMffa4XWIcZH7YDpuZT2+wtqJkk0proTk6ZuNNX+KCeNvFFOTFXyogtTlfwqzK
8ucBSlWDAll+huFGCOwxaIwjFEiPhZMpqpkZODI3hTNj6xx7qVl4dsRAaWBFqzqq8668dRHk7snr
ypTfrmBBfxa1ZIpv+LP9aEbaxsjtQ5qMkQEV71EeUkcQ9AE4I8EDgmDblbKIrn8FIjvWXpaabRrK
fQg5pwje55qtMcm+x2r/rOapTR0/2xK7lKvm02Dp0vqgvqSV196xHckK430n+aQfMbL6obvkrfSV
WnPz66GenyzBX9neDp+tkfQhhs2dXyq3RtX4YqEcKFnyiKTtyALEZy8LrWwIbUo76M8gkSH0TBCw
aQgCmFMK05T54kQmDPyczGyI5GjvRgDC16D/J6jBlNoDoagmaCdJ+Vp/0bV2Tgjmgy5iF4bfI/LR
4MgY6ubYQ4N6MI8Sc0x1UWxnmLMT4pTfAzKUeyD1gzAHJkWC01XXi/687LvhgCiyZVhXo9jAOzIc
zWzJVR2kVoWZLPSdjj0myQpiI8aRU7L5cWcMrQQCVa5ONzttaYmicqukBcXRU7ZIeXEF2VMl/is5
oGyG9F/lPD6b7lq4Etd1jPLpAjmmX8UO3UHqD0UBOGIG9a3Rwz29ULRJdR66bcJbaZ7aDo1osYGa
3gVvI8eqCrGsgKE209Dy3Jo4BS8G1srq1BHvWheydWNwfQZAU1Hibh7fRDVnXawzLa1oXGjjvp1P
2MTb1+C4T2LpHGEVATIeLMsarLxS+TkjgETO0HWHci7sg8jMBabElbH+p37qovSbMIvu09YJHz3j
0SO6leo7szEwYrPOfxTaBZq1h8DUqvdjKOkM/al9qts6TrcnnnygJ9YIoJieGuGaubgEy8I3VtER
xEDoAGxe/SSUyvHyk0aX0Hj2IwsDT0zDLnhR4qGXQb7WPpegy/xg/OWBhVD69/JPLPIsG+KaMRoJ
8ABYmB53fKbd5D18hYE5pGhEIadIWEtfwQfjaBT5mV48p83r+MHK5/JCQrvoDMkyXAJwt04NRIHA
EefXEnlCkj/YeoF0j97sKYZ1NCiQo4hmz9VuPUn3i4ssIjpJlcKXyuyHLC9C52yxtg515bJllGLH
oVCHMgArh+k4sGf4bFfqM39b97B+6MBXkEdvpO7InQhfXbq62rGEZkAghQFRVzTl2g3NVIo7fcTA
vvPFfnSdMHMnqJMDxRCY4mGGaPQpBsaq0Wdbz4H92ogTbMSi6mKsklSBdE/ghT4M0dxzJr85Uuff
ftfANkM/ZhLrfiFCw00538e7q/jya74qWeyeOd6tNJ+wteKlZMfbdbsLU9bIo7+1Gi4XbHTZ0WSv
GHbx2QcSCk58c4Bl9fxdczeD73FBhDKq6831glhoQknxD8ujH0sdozxVNpKD6uRmpaE2mcpY5WvW
YMbKuezZGQ9F64hptVfSqowXuUhuuTfIjpJSvpn+CsX3tFqwgl6u9EY7JjYguS6a+M9RIlcKqWLW
YQs0HnWetQ55XqiROzlPDsS8nnon7dn/w7JQv4fFTMo8RQRJYdYIa7BMo/+shFjrRW2PwuSQ/1QK
55Ne7D2qTrqlC4RVz+YWz26/rV2hCq1deuQXMrTBOWcuD2fPJKJ/z5aL4NYNSItlZYiOw7ms++L7
1lLm2vsSe5jjuBwqttcxbmAWXKh8bnJH2+oi46ynthqBhYgmhgyVjk5SyjtdZDgdOLBxIDxIvI7G
UlGsUT7+y1IyDod3uCpI5WDeVEkrrQxVsb4o9D6VS0SRLuQ1VKzRKDAmXZinYaknNIVaXPfSV9Nw
/7bUQmpsYx2/lAa9mYP2KxAJLD75GH9vdaKou15jKM9mDQ2JsYMWMDga+1n5SLnzrUUy5WmX/OF6
TMoqmhJiNeGMAfM1npPfREPPLBEeclhE+d7UqHZgl/3G5mPTkFdv/y1GVFAkCMDpqL64sq/ZAVz8
u3vlJVtpkn3QvXJvGisTv37HYJR3Yi3yS322F0fdsWVJGZyNs0OFeoUSE2B8hGJiMruCBh0fDDz/
+wt2yvWmLSvKryvkNCj4iKC0jUwxyXNt4/gwpbq5e2V/44IAJ6Ax9fL8uAqk2pWmcZkSUd5iAvib
N9gYsGhUb2FyqBmYn9OCIasVz52ISZcLauO4B70hZwaO3YnPYBaDq/nuI1JCAkj8pc4cRC63HRDt
5ff1/ehUKDGDcUaU9IKHHvLRY0SdbqiABCS5rb6QwDr1ktx5irqiWJERAPnLDffrd0An3HPoMTF0
AfpxYa5bWSQsgvLcbynEw6Tyd4mO2lD7NAIgLE42mMh6/dyZ+6fcSbCK7gWWpPUH5Kv+4utHFH3s
XSMuY5KN9XDyZrOMweX5MvX/ntUiwx5+Sq4SYnl7mGDvzGvcMJGFBv5mJb2eR6yZLKbbHgthIS4j
pQhfvrfDN648iCNbbDdH0RmQYzMlH10OY5vEoeDXGWlCxJ9w0Y0S32X2BgGhGCnwUEqaKIFyPtPF
YxJj2SIB28i8CAJZm94pCv4LL36CWKSdRJCgWzVslnNMAkvlIWz650YNt4809p3TioUN8lpceZ0V
yDxnb2+dUMpjcFc9bLqlr1z2qfLyQxwDpSoizoBKwYKIpVkK0Vm+FYtWwP2kdDRgyMyVDVs4kSUo
8GClTUF1gr6iwpOUnwEyprG3ze209/pXiOXq7ZAl6w5q4asgHo5grT8kEfZZivRA9WkjoW7HudwH
+8GwyChaMPIJBvWE3ruM2tI4yFJl93hsXhTBs6HdQyrni2tB9UvIAjAvyvo214RPth8BKnPy+xMf
tHcLZIe7tSA65ExdRUBz1XHFYBPTlLocHS2kcKVSFlI3t55TjPzeRtjKpuFvaiGeyAzIfhkqZ/xs
yNPehtTBsvC0n2ik6+j/AaFrbNscLu+kpMqa8SABZEUvh92AYqk8WS90sZrOuGP2WuFKaG8JrdE9
3M1wf5WKAF4pG9CsqLgzFIrBqNFGb33UX/NdE1Q0NDcMbX1zI20e34in9IxCM0rywqmb82EQsAKP
JtzVktWlcFgk6PEHHnEBlOcPkLaTMBClzkp98H5mhc0IGvK41my7AZYt8EILNzjelI0iqyfOrem8
DUpVCioDk6ji+/s1aTh6ZSQ166fuaehWmHxzmHMYtGJF96bVcgXH1AZfWaM9BP8HbYf7svVdOk2K
o2OTO4+w18bFMlyTZbET2KP2Va2WO7tyvRkw6+f6jcTFUyFl8lT3IIE0zaF6BN5Ygk7xPkNqe0wk
NkNeF/hZ+pZ5oLqCfNRrZytas23hmSLf9Lf/gGHFo64im6ytgSS6x66Y77xeXgwZN+rDXUSD5hRw
RRFZSUU5W5fmC3IvShk8smsEUvMLj9cmhETZSMI/njcUQvkXmUJ/3b+IfoP05dmVO/aQamkKUQQT
zKSXs6pi+tyoTnDqQ694g/6xzfUkfxM/fr16cqU3OZC4wuao1+F7wAXjK3UuxnSw1EQwQYAFW6Hl
RGA3bpwU0G0HqeFLBdprv/PjrJq64oKYkLErAaeIhVgs6a1jeOBaWGzks7FnNjKZ/p23X8zwqoG5
mLimVNSLvLP1ckC1qhrTXVr8pKd3lKPnwxaUu9x+uojuxiznrLpLbRGx60ENuu4E0p8rCNKo9/i8
Dik1mD7/PLG3zD/u9bqQwDETZn4dzxDH7r+nEx4gZnndpw63nXGK3kK97HkJLjhjGWq7IRl4NoTK
21zNLd3fV0absPjSert/lyiB4kfPSMxnyWjg5vJyuweXtA3nClN9kOLtYkOMfMuKeYTXLV48uy9B
Wqnr/LNbV91bazGmrL+XhgZ20lRwGDIGlT+tblyr4uXcJ8PZVunGOlHwSJVZr31CxFmJXdzIQ21u
uq1jBIsaKZ0+orXtIXZqg0vYgKWuGrVtktHifD7bvwQCIHlTWgWJcFAu91qZ1wMAhZ7oxmNsg5Fz
uyMA0RAVzOz/wVHFm+5wmJiVyellURORqm+7q/JGbBR/YRTXGbch1tn6g2gXMlJq0aD7rAhMzLBW
VcQUE9+LpGr/ONoLBd6jltOwXcFjvbBzE5gkIoLsyArz7suDqrD4KwmeU2yXADtBi844vELV+8Ej
3RDwfu/E1qRmHR8jFXgGEpsoetv1uwgsKz0qsmCKMtRAFMsDvRXhG573KXJQ+yGi7n751CObICeK
kdX1/DfmULETYJeJuBuqGeYJUrH2zd3BLxenomtive7O7kHw5346OvSSwZ1hduxVlp1U5hqkt7mo
6KuKGruO8Sd9yp2PLdd44OToTVHQ39DlGfpC0Ta3YiLz6vYqFsjc4KadDywM/M/+OJU3olA0KALR
mD+iyXyAvEKvZ1SRh+Qv2oRNy6LWsfTD9+cfkMoWOfFF1+GVSyQgELibIrbwBwrbXKNanvmi5o+e
3DK8A84zSQxtUr8R+IpMwjVNBazYKhcQYwdrjzohMW83NwMYpX+DM3ooKUki/tCVwZ54m8WTio/7
OVrqFtqVnk9YsrzfdpA8mc2YiDoNCkZqm4WLsoBGfS6zYecRgcXsE5cDWjS36vtH/Oz6au7vpHPa
33K6VJjZuyTIk5/UPT7AQ/1J47QOSxx6F3pySadKnM4Yn7zewhKl1JEaAXRCWixTI5JFF2HJucDO
XRt+G2sCxhSlgc2Yx1Dp7bKR1yerHdr1fCQB3KyapkKGb8mt8ROFo9cq2b5q58M3u78FmPjo7mW4
5pKqMm2dVjKSzhVg8yz/CPvlMmWArJZDuDSrg2KN/3WFo4iTmRqt2TmfTKjD46MtY/ARk7/qoOkv
qXmeeGtNeoLsk1gWjJaaoFYhBUSXrF53xCvMVkqKMATnCLvhb1g4rfxbDsjV19JgZ4wh7TAkGz6z
igSFIflrSKFyrrMMDDYuL9JlVpP5ZzytbwkrAEujC1u/IASFX0YzlFK0QBHRiDZLW6zETpkzIAom
3G2ECn+pLt8NhbcGH7dthtfWqUCKIfscW8XNszk8ejjXMwY/r2RMQMfVu7ghl6o/yOdoQNgzC08Q
pKqBkQnZa+7TUFr2A6Yvkj10tkeOV0g2osH7vQ4iqzpydl36h20i9Be6ytQJ9hi1oKe/fWCzJPqQ
MLnYLcA7NBwPlvn6Cqk4B6U/NME/Vz9OzS/kv04x5VdBqn84eogEUCdT4TMrvxLnMW+wYVtAlF4u
SNotJWNIN8RcIpw472BC21ulcV3TMjeLHOCXC+mWFFhk0yaX/KZk+e1FjgXfUMfLZG/hHsuvRESF
tIxjqWApf8vAeaOkhH55An1+qFaYDtMQ+tVUQSxPCTeuaIiAgeR7LYENpIKGGYFVPspDduzZX8RX
P0woN7eqn1I9dboJUwO8v4kUVYmHUnl01R4YW4Zu+J16J66MswXKtLtOKFMpD7S1RHxgrLPPUDoz
S+vqnfxYH/QtRCtCcdIchZSwIvN7Wx5u68IiJ0rRfG07TxgUKxn9hFhxm5cdsDUJw6YIzusr4KBC
XqxkkgmuuFeGtQA9h9Jydh03IDn0+e2G0QvLA8jmdJVn7xevOYrAxpDz6yIB5HrWgKyGJRj79mB2
/6QTPzgPJZHlIsG07tkZbQmJ2XlzkGScxnDLh+MNGiNKcphg/9gzR8QQcBXTPgwI12qee6tKFJov
WggEADCZ8EGWlYId+yfwbOYy7/KPWBHWeXt4FX99Lae7Qpy/WHwnQfElj93ojOsKZnxSfNISd1OS
QVXsjWNaA/wkZGl69IHL7/ark/SdxdDKUQvqk7yEZUN+ekBXad+cGR/ZVluMFIbQVVXk60h1lZ+k
ddu27YNOhv/V6nr8UeDo5owSjdaYFDjvwuJMYY46Vq+oHuef6Rn5E8zBcDoR1Undznlr4MjguB0q
H30jkirR2HHzhHh9eZirTy8sX1Lgup3iO1I5ZQpxYCMnxojXv/DWzn/EWXR03sAAbfK0etS20YqB
Sdf3G4EKKFnLHnYMeS/JxDEvoTHSrk/6FxGJhl/xNBwzLt4kCBgursPLsgE7cbdytEBKevyL9YQu
bVYIrsvF/W9GM7afI6Ut5+tgzkJ3rRWgNfS5N1qyU9d5rHHhP4a8ApLPxoxahCS0IccZlFG1Rgks
1/EGsvrzdiq5Q8gtHs76sU7Iic08jM7YeexxTmqFWkUVoe1wPfC2FgtV+JmoUGiBErZw4zSFdbvL
NGF3an16Uha93Xte2HIj9WAYSvlxKqFlZf9+B112xE2ud9rOc+qXk72kXx7pe8etgLIZVDiQ4652
9tlQUpDp/3oP9IaO6TCuchbCkzewTcWVYTe+uY6YmRrKiOBMsab7tQuO1tEtsWWD1PxYaHulzslQ
vQs7eojhftq2plmn3jDZ5qfdbbvfNJG/Zb6YL7W1fQoa4cKiZbZDFBg5PvTlTtxgrFOQV0fNC9TW
VsPHozJbp173obIejH+IvWTYiddaA6QoMBQzqLhaFnaGOPU4TXvInmeN/ZhrxL+XMIbb1mUifiXw
b40fSkphJGoMRbwJRKsmIWSrfPoUjAWxejNKmMmWgGj6J2Ei/phSg/m9uuZDJM6AOaiTTN4+qBgE
0+RM7D3dF+DYEVujarsaflvcAceBYYR3Fs8gmvY0KhlsUejaIRQ6z0Y3gcdoKLQx5DT63a3OY43h
MJoTeFaPTfiA4gTQNvqN69ISZKLwOBgcrKPj4yCe97T1G2dx7aMu8XNAcMOpy6Y6PnnzRtkALahj
Wx3zxA0qD9giYTquXX1hFMmdDb9iDvLAIXGJU+EAGe8eDMKwlaJs/FJfSJfdfqDa23Su8TvMCGTb
acyh3pIFnRwOtYSjAvu91gGFkltUOM8HgCUmP37YGMz4xctGmY7x4hBkaJuu1s3L0j9k+5aKauQy
UZZ7MBWAo5lUBkvEmyJLThLgJkFiVmnF4IBzqCEY9sOpuWazUTTkUlEue1MJtnCJ9sLV0vJjyl1O
Fe5O7jYRGrRjfJFa1q4Uz/nOMdzYephxDWmo6Pu64XNVPOtXPKByQeiPtzQS4mWLTHK6AfMS1SBF
pQcVjO4JLNEZNcCkOiAFwH3CEITJh0YtUMQW2z/16fqV2gm35CPR/SJ5+5Eff2huZO8XMm+GTBHq
2eS2V3kKzqwZ5ZjifTMTtDvKpsZCVmkbVcHxTAZgMnlps8rMwyGwUblcdtl89rCFNma2mVbKsVZT
5A9K9mYMBgL4y24RbYjnS7wHqSQqA6WqIUMCZAoUzsV3vpRUijJmnofTeQ2JQ4IzYuJxwmm+oI06
8bLxD+ccXeH487SlWy5hzhq7kORZvmeq9i7DN2LwMGipu5FuO3JZZ2I2FUny/S9dsh6bB1VjNKNF
dEPzhPLLugM2GJNgFa4uc6fov5b+NAjDNdOc/bI60J4gjqfNFvIlFXqewc+d0ORg7r2iuBH7mkEK
NU5yt+mLeyStxKi0xVRO5JuKCBGMBRZNhDc8ih6iSWl8FXsJGmnswug97pCfrXNl7pzOJi/iJb74
E5NRM9WDmsvfH3CPDGjPFvRgUFpkptj9x4AlJ9LstPAt5Xcf0fpLkdHfFcMejowqR3aTvO7QsGKW
hpnAeFNK7hGODOlmb+bZ0ZHDRx1yBkpI8SGnOdrgUqLvzzgsBRigtLzZ5zp79PNq0QTL4RCdVd20
wnLwgbJMaz58WnTK+oyUvTBsEVUn7OOX0jU+qNyvIcZY69IpukpF4xFfi2H+0RRTc94KRHdg1rmy
BmyFjjFNaISCbNOunYqWjG1dIIQKFrCbXgNfHYudeNm2WbRW6u3MlhXTS0wd78dx8N69LnpMfa2e
t0w061hxmI9ugshCzJPtNqURn0clOPqPLMlJkRk/x6TkoKbrw3Ue5Ei/w9BblyMU/MRBLS1vaWlY
BVV5cf6fNrjVIQbtkNTW+snalkn3/MwA+/JNhHo9Ykm2nwmclhZ74DLBVkKWvkujpTtbugqKBC6b
T0M1bqIxDHYgekzTVK+k/ztkIv7ofG5mi9MDPAeCBzLwlPmo8b7AUZ8n2jV/NfLfiL3DMWyj2bBL
y2r2vfsVlhmmxLVw0Yw1T04k16jQtWVPfyfZGmOpFpi7feBvgxCUEGwgCmXXWPPmK/RrbGUVfxjn
1ituyqdsK+cxbLo3RkXO6QqA9Z79ihxUcINxgcV61tRsIJ9zdmoKcOgmLxiaoaoZlOdzwWWxVkEN
sQSardYGQNbcoo6mSzyst7XMOAHBRLoAQ/EGb1xCpc0Qnfd6aj27jJnb1d7UM0kicFp2LbEado3B
OmB50/xL3Wex7xDBKJgg16W/rxPxBp5CAY1Ct6+JfIbdfv6o1nXRpMP/pLeRS+w0R65hKVRvrgV3
48aaYtqIvVH79XqdN/P//7D4dOa9ujRnPfK+CEX1+oUhlTN+2mv7PzLwrpkRJBmSG5UueZDqAc3d
kPro2X9+m4sut1gTthBwpGQuxrOfRk1hu1W3e2ovmMwNMRkJcYafIfc2lVtGAcfpg3XRbLxgjiVt
vhVnGDq9dufqvtTw3FDH1dGAR7eq8g7NcRJdAfy1Tnzp5uKqo07PHV64Vxg+uZB9Nhi55pAyU+gv
RD4yVOZqOZuQRnlFK6DYl9shWQGXLS9q3rBd0ObuT8SYevuFGJGNGj40HIhU2xJ8ol0r1pdunWkq
uwrAv5C3uwX0z/ntJt2vMQsEu1YOcOvFqX/A0micEG+68SHdKLoQOClaifF6VhBRZntDU2g88Nbq
eyq8WdCyIE8DU2HsH0Lbh91BMIOHtNzA9HSg1mHSdc3ItF088+ZicbO4mi15C2kbmf6slqf+v3EX
n/jm7jOiRut0mYKu10c3SQkVxq6uHXoB2959mcI7iX4JEiVn5DuRBvZxTVuS6K17WLM5cQmFEpf+
JVB0nfsIjtWDkvn4SP8R2z5fC6c7U6drarbKERv2F/ng6on1pvhw5traUcDDpmihBm8WsNpqJ6bx
xVOrmQ0/1F+NQf3SXew7+NeKFzCQIqqo7ZcZ/D0XDPUcd/lvv0WDpHedZ4+aUmTHLyHvwXg2WwF8
D5Z23cddCwTXjoXvMLfG2dnXewk5pfx/jlUHJo/PE6NLDTu6gJ6JndLWRjG/jRS6m6/JG89QAdBe
+Fm6ZCzIIwEJPr4dR+HXOiA3yIBOigAoSIHHx6JsUoJ7BzdFfCxy+QY+ay25OBIzmrGVFx4IRP0t
/x8z6Cq7aYDdPsQ2Chg+k2OPkJL1QlnF7Dk6WTqZ8aH6L7PfNaBU2bocc4WgNP3QWtTmsYTdyFUP
g7DU0t/+yh3X7OZtYHj8VC47Fr1ai28aVMrmx3Wie7QTsmUonDmTqtbhIbd63BtECZANLpqc5PyH
gzCosC1B2TPBVVMdpsNQtAuQMBCtru4cAu8F7qdN0AMFDs3xGmRntFZHbIN65dTuyBe5xSwFly7C
yu+9S3VpgJ6bzvajhQA4BYiIL3b8yQ23hVm6e1dy4lGvBPYlXs6pzi1nvUpnCUugJ1GQP9ZKY8mq
Ki/1tjuCB1itP5sLUKV9llhHlTsqZDqiwZ2CCDmNOIwuTI4Udaj0R3DaxWXZRPk03H5GIXTByAeH
EVC0iIYZiT+VfwYmVDtD2E+PuFW5oEeWV6zs9M1IFutNZGF0bWMnSOppDuLB5hANdnwQpodsbFbp
QVvD5jn2sqvHXVDJgXL4xxotmI5VE3qAqfOE2XMmqJ5eN6yAyBxIHatTfR5qvHr3G0C2wQ/QVNjw
fa1hV1wlLVodNrEnbpQ4+2szuhksi1zi4QHLLPe6v7zJqLFZR/TTF+eiWOW3dqfwXkXTJlvei86L
jsVNk2sBcQ1xnoKDcqQMd7SFGEgSWdMrqtE59R7XkefEEZbkdfNUDONeTQbMk2wOTNM2q6rKv0Hy
no3Hn2Y32NwsFXP1huFpw6eBy5qxkJt8B7aP5dGwQMb2bEDdYown/GXZZyYDjjz7mmCpAg70EM2a
ioxAH+4BpU86Pqj7UvG1EOfTDX4J+g0HoYBEVne+v51Wq9mmDiI+AaCAdwIPb78feRAW1AKzmZve
dzW0Sn7p3UkqpAZMIin9NTReCgFIEhbMW6p52OCfSqdGX0c3zPeGHkDXYt5n2e8NPsdSx2H5RSrn
5tTA9eEgTXcuYA8CEkz/2//1V2tDgJ33fO4JAqcBKA2HARlqFRX1GGIJgTj0ehCVYjlkoeFEwQjG
Wd8XVUBNwjKFRomElh8+cg4srZPPRHKMvbvzHGTa6LA5jlpTKp1MsdCoEq4UrvWFvqGFxprc5fdP
u3GcoHUCUR5mYs+CvVAFE4/C9f8XAnQLgerJgiu4QYVYVhSsFe114OMH2nxFiybKIiOlHraCvXC6
tTysONqK/+EpIMLBAorHweOqj5T6KsIR1GOQRgbjMUFpAZ/oOcNc3YqSgArZdepWzIUskXFzuMb9
AoIJUu2zxtnuROJRcn8bfmZjM0S6kCKpV2E1dk7L4XGdmlU8ImsE78QURkovGuaBJGbV+N+DSqhu
9UTa9mXf0IhhrhXRSpBim5oo84z4K4vqEAeRPuRLy1tiA4IuVsLfve/obOoYNpH1rlJLMDERHyOb
9bItUgIJLW62Lez2tPIorVonX43FbNCnS5b5siDuhIAzKeoCB7Bimq2J6p8KXqFuEhlhwzgBOEkj
8HyH082aOXfW8dwVKPz/3xDdxyoYA5+7m5TkxvzyhI/v9UvNqJzC+mNA9Cvf4+c+q7VvvHdl88Vn
miVeDt0tWojz/K7lb738N4HF1E/+qZUB5spp1zjF3IWc4MASnOQAvUUZ1s2guu8C1AuhAByrRuQg
5G3v1mekYV5xsV4/cVV561+Fd6efTLwPDcsrkocEgdjLSxRxmuw2rlcIhn87YSGQCt58cHeVgrte
HisEt0IYbKfmG8mQMYCvnkVTPrI9FDqjmF/pJoHpAMQB/Q8ulCnziq39lAQUnH8SqVhdi8XF0AmK
rgPW4fPOGNr/nu+K2IdWi/lD+BeJK686H901Ac3l7D5tCVbW/VkuwlUIztpKk8QsjkPM8hFm2dFf
aUJcMkMisyU/ZqujZHAsBdDy914tZ0KCznNVflGRYdI4jTSLbA34lyy1EQLHD0X+3xkp5ViWYF4X
5tkylIcstlq9HHbN9tKZOqPs4r5f+29NhOE3iY99WVlkZeiS2JlDTe8PkZLjDemLV9zaJwbu6+fu
oajYFl5r3gBEZpAgJ+3ZW2s7DlOusl4js+L5zZqJCYwrq7qxqqvt3SPu3vd6N5IPsXjSTDm42Wbc
86zJW5jxtsyRAybXwZEN3eiGduR6QzAYNFnnBAhYXvv1r9Bt0xVG6S7y8k87/cm80m9FvUgSzITi
g0/NWZijEEUneamXKVlBF3XytgdeAWl+KyNlUQR5O9EqF465uRExmsSWyiJ24FaJNdpPwmNZZk1K
8pnPu1K/3K1xTkGjmWh7a28WNukNmFPgNmAyGdkjMdg6RLf//YTsnQ6IsY2YpkijEfXWUGP4Jka4
0XRB7WCrbTZY+b7bUsSYq3ZkwjAJILBlwW0GmCoT3i+DmienO+7K9X5QMrSr4L2sfsvA4RnhjST/
uzegoe504d1ssXmodnkrOaUuGZZMfZCKnpZUuj3bGGqFk8NaaAhQMqWdY63Xd3aNWTS9+mUpZqul
HPLE/X3+UBq6BJsPAiKSjtsNhsYnOiG4wArh/EdZn5Qo+PR0srQ1cYizIRzzKZIrrKY7ZcxR1HuW
fjtsVjTMgFZx3p9W3FyQsytnAL0nT2R7MmQydztVgwE2Vsw5zoP8RLGjJeAICjXyrBrfS8xLo00/
zA9Ndxt6zQFnETRM3nAh70la6DUKxw2BlSwYqv8SQDvyR6FAuE47Ynj37ZZueuFjgs/oEjs05vk1
0FqQi/2x5c16lMZYWvNvoAVWwthKA/uGHw3dtgRmGBx8KwYnVJduSz8m+n+H1WJ8oq3yggpu6WcK
jCDoYG3P/xmKJ4EyGJ21juGgRrbQdhH3bPJDXk9MKkKZ/ozz4vpk6zMna5ABYaCnpwMXIoq1zVJU
2t8RTLv1j61Y+o5H7BhBiT4KCGn3Y21jAjhpbMISAo5PaO9Q72OMKE8qZWRAN9OXLmz61/aOZ4DR
VSXkVXv+tuCrFHkNDEknTkim8aNHK+lf76p3s386G3H3rFuLMm00vZvMCYmuEF8bZSjfUWAQyT5E
o6PvZtvRQ/It6a8JjGr/+9S+tnYwn36BILFIWQzYQ1gDWGD+AVIKU0p8ahYqv14bg11BIYZae6G/
WDbpJJZdxaVoUP/v5VV4wUfOm5cB4kAXAilEVB4L1FdH7IQU2iimYXv8liOqOnv/4XPvsq5Nslmu
T1LeZusPZDl19YIA9rnos886WVmgwTWS/ipy+LHWs5Wr7jQGrYSloAjUSM3Rx2UrgGOWEW5QEwKl
lcjTz0hgmsWgiPBGkT1x1c7g9KdkTNCGxs7r3p0rpApbrWNv7Me73iyqCmgi8IMbnIlMmswMoDuA
n9tpzVyQnfWVKoy54icBGjHJA2HNtr11hY90LOPgqAvn4xgtg+G/+fTtnU7hpuIN4Zd+OvNHQh+M
e2SkLO2OF76PZG1KtnMaOPLFPqHYxiJE/y5kz47PnOSCOMJwXm5D52Fte6fvhvXFMYryveppzms4
CSKGp/l9M5U0ehgGqa1GmjaRF/YPd/0G9b9jFJXVFT8LHDsJV0kzCS1noo3YsJE+V2AKqfCytrql
I4KdXvs/mfkJWTTDsG9aaBu8HBsTnOK8FydtbyjYzDLalx9OerAMU97ioE8FVfHqY7AY7doApQYn
Mc6tAnhUpW5eeU5KKC4RcqjLyfbNtOilx/AvC8cieX813nj59oTNFiqqtsZXFd8KiJaDQwBucSxk
SNw6k6Vvs8r/xGtD2FEIsDAHaEOwShcwwSJzYcMVsLJ6PRgwYLXk2CwUGhywmLpBsg5AqBpAbg4v
LidTqhfvwKUrAbit6KgnOqaRxY1MNKI0vLPwulz0KjCVh/0Xr6G6hRnpPsqgX2BBL9d2Zo3rWQVY
r3LmY5VvWuoW8Q3amzCqag2nOdi3qrzjZnfW6/Iy4jNPE1GqiDpflOahOA+mkAa+9fJGmbQoDWaV
xgipHBk6elXmQQYgp2QZ6R9IW+Ls63K+0w+EpBrax996OWWzBqBzDcjS0d4B7STakiCQpqewHnj9
cM1xPFmPVZ/h9FcJmF8dyAgCtnO8acWvn/HBCh39kcDoi2BpADHEpzWS30s+wgVEA/p2A4VefCT6
V5S6UC0K/I3G2W+j1ZQWovVv1mz8U8WB9p6zDjRu1U52EWP+ZzyF1G7qdYZAsLsJ+dRNSvQu8+dv
H+ftCx4ZX5svriVnk3cMa1bKU4hQBPC5rJGMaGCcBVSv7YTleN+OoHGEtCfCqs9P5fX3dnsPSfd4
ELORYkBa8xr9ri03XJ2UNdcKl5g2A9Lp9wrC5ebbrMEeg2S/OrOvUS3u1hlsh8q80nX7VsLXjLKD
XJ1/m5oqU/UfBC/lYRIqvSfg/AsIu69WMA/Ed3z5x5LfDE/jfGcJtMNKFV2UUP6CWiG9jW5TaaEl
WyHQzmy3c2MfgJppXhO43NfvjMhj4MMuZ1GH1Q5zvOaND85Sdhzl4r7lJy7RsAsGamnbfML0qd9N
abGiONOBNlUJrdtUjWkJMbyEnJcLB6LPnkacFhStiG8sEIUhR9E9nNGFAtIrJwKmpgThZg7yTBmv
3HR12W+nzY3IQEbmkWgTFpA3kgjP20EPE7cZYsWAZ3r8EV/BDnGmAGxGR0Qolsi2mGHXP1zn1pdR
oSjGSNbO1cgMPP6QHU2DvbOs5/aZgaqISlZqHMrHHMLfBECIpGJCqGiNnBQR01n7wHD4q+W5vCQH
WzAFiTUBmNuU2MaJ69FW6c1huRX7MdZrtd6aOC4WvCN5xRyUvSWR3aVQq+Z2i2dQMQ4CzntsrLHz
8Qh0ijc0NA7BvlthbmR6sntudQ3+wNlVQuh2LkO2R37UI5+MHrge/PViqfBgGZ65ingOnxmS2PEQ
hoxbzqVn0ibVgSqLielJ87m472A7PItsFiMVnjipk7DEtjq5aPvHudmLRFSzaBN+G0okCEwPlHed
yYhbIDGs9Q2Dx+OVULYHpSsv3uwnYTmhwiDPxwIQn7C4E1NplmQPPaG4+F5aDamm98LzENXcK1Nh
GrPxAQoUcb3jSTufBDztBnrjlVg1JdEVJPlhBBZxgKyjLwMxivx0nJ9AKVTXfxK/lt+PrtHkLPN5
iGSeR+ubdws5ZRRHZweLLiY8RX2C+K1CYTR6ay9B6U28SxTUFZJI++U+BKGJ6NamPjotI7kt1+JJ
BRW4bOZVMNoFSV+72u3fah60uBdGbwbi8207iCYXwY5SFSekaURPF42OLoyyzU3M9YFiplDJQorc
ikiL7Ma7pHond+gbnEZVA8D8iavd3VuQx0B9ext4q40CeU/iTncP5kkVb6Y6WvVUpG/z32pi1zm4
GKwcW2an69PhOD+mUTFjjYpa1U1Rfv840ZvuJ3dtrR/5FCQQAscerVyKPf2j7DcgPyR0ZhCKrFDk
z28MAwohphrau4RULCaO/Hv2ss6zQQdyav1BGlxPseRIQfSC+egjOr6PMuutUgdl4rBakXAnQ0hE
I4VuMntj2/f+7CNj2hZ7SO3wZacG20aNvXF5cKlmx80rIB9DU8tB/A7IxqwDphKIwOHCKz6sX8Hh
Camae+c8nOYUyuoS53B2zxH75f3fWihvRQrwaKVKthla8jdJODXvS/Y+ezSur6QlWTeFwK+eSiNK
Qpqm5caaDzosPxdoYhuP27IY33PWvVCgjNI6J2tgQU9YT2SyUc7pO/jp/4alQlaa7L4wQ4wsuKug
zG5IrVd/0V46lKS0u8zgeImhIzEo1TT/yzGpgzIffIIODjLL7a8pRBycGDQV6kOd/v/tM3Y4A0qa
Rr4CJy6mp/ETWMQTt5QMOvh1BEn7xzUXDUv1gvoG6zm2Y9xbr8ISw9amGBxZBwlTCqvfQxHF9mln
h4oGc9WmUgtJexB4QrAAl6Os5EKCkYXYCJi0LYP4zOdIKWXimZFmV0qhFpf66BvYCIOzOCdxWHbB
cseVDLy/I12iLR+G/e9ILNM5QkWDra/um8hWZ6nmJuUphEmaWyeUdkDbQJw8+UrGpgvUjgWT3FR7
xu9mDE12+uFEoz6Z9Exn81d3v6xC9SlAadqEKjym3Pruc4MHMQzZlP49w05uvLlm+cA52rLsg02T
7z4ZAjekMKRw+ejrnxYTo+EpUaT5IxFJny2gFuUNfRzD1q8siVXrenFbtPGhOmKdhoe5yLACatjs
9TjSVfUD0tavQwRtv5JRo69V2SQ8aq1YkA0BnVQXxR2lLU3S5y6d4+dOUuA31Gu8eYf3zX1f28rz
JP6DT6OBcxbzxLdUtO4tfOW8e9Ge+jJLGBXC/FQ08GIBfjnq5LAUd1GNtVhxYZT2EAGEPY0pMNvM
HJl0dhDtFPcrPRRSZ48jZt6+xw4vjlk6aDTAFtYAvZ1DBdBFPYRfvoYwkjI96BwIwmRkuE0qhmA3
qDhppBfU0cZmEPTqDQPNwmSYp/X38r6vrTK1dMcxPQYpPs1AydesubSh3g77tyqwO8JiT14fboH+
jTS8Eu6VQXkmbsUCJaBfWdKErIDh3nBivvUidY4zNNfgxVTApWCBN9nwJHM7ymQGQVp+u5T8VQyK
Va/dk8B0Q4LQD+uN2lDPVqO69C+edUrXWQ8Cm/XbcW8FSU6K4bF563I+0GFdqoGLDpI4rQ5LgnrE
4erL4tHR/4YgXcVpDPMR4p6casmEa+vB6J+O35jfFOAQYcF5V70KuFs5QBYRxYG61WZdn2d6vP84
FdKfwQbP+q4AIxDYGmMCfLgI9NTA2zU5qXjPm+vDdXWPpz2An3OF3zh/oGMWBwjLdt0hfwifg1xx
4+J+RTPVs7PZV317i4JgbqJkNl+dDcZi5CVLEnynkOHP3xrrapvml15nApVks9ghJfH4shyFqiKH
ITNlnGXnKnvGmRXKG3XVRt4tiP0YPs1HwhTIdcWcYuqJco+ROeVgyjkiCO0g+3kBTlDBTG4Kz9xr
oYzKJ9tg7YJEXnADXZAoy6EowvUVnKDqlnBpgIHqQEyW5e8bBQGZJTFuGswlZL+gt9lWx0PT8JRX
Ey6Gwlx2KTcdDHNs9I3FtZEXyTuFpahFOlfRYF45lpT9U8CmIrzqTrQ5IEyTUaaoDFcDjweT/+27
YoEIx/N9f4hF+b+cgc4vML/9IsdIYqHxo8nFyeLWrgtXwsHE9D2uSQyG5sJZvRF671BJEZ0K2k/R
BfmSe/DA9sp7IfGniptjkVxDXookmIIAtkX4lVzqw3NuTDT3LtN9ipyImB47SUom03i5gYDRnvGw
he0JuWfkmhMQwWliujfEvWpayRWpJ4ur0qqvavejtSGBrysm/FV9raCZWzonb66oeCHTKNQcMnuh
Im8ZPHgo3xS/PmDD5n5/CPdozw0qmYTp6ZUEkHODsn7YPC3SWK5U/RAwIg7OMBZfw4ZuAMrA+PHV
fhvJIM8zD4tMiRnXrQ41mMkOB6BbJkQBIiivX4DPYAQ3vHds5j9vfcosNni7PNXVUW3QYr+3kmoT
rPtEpZ0Ba0ggSDUxH+neu85dRGTwgF0CysRPnq1E7I0PnkiDLv6ntaoc/Hfu5O0iVUsilw5kydzo
y65FdI38TdFBSsV82xZo/kEZdDtBMZD+Kx2cj8qBiEOcvNv08XJoaADQsGbNjN2+MeWtKRH5v9w+
DZE8wOlKo3Dk2BF9IY8izXFI/D1ibjb+xm3sei+YDtzRNVIz/IEHwHJCmAr5K3DjRVy5bs6qc7pG
Clyow0W7CrKWuwIuzZFf1VhLC4CNWFAUqrNWob3gDNcBlq27Oz2Verr+FDKQZOS4pL8D8mmu7H+T
0BGKFVIkZO4Y9+QwXSBoc312Nby7WFecbk71TMl/vpUBeQziybnyCyTBn1zEZ52pwLcsZQOUoyun
2M+PiW+6o2b79l0I04vrzCDHyLLjAhgjc2hUOLCd8xb6hCFfSvL3dipb6naPe3NcOqDzqLNEcq51
5AOa5R6FDNOxCxP7aIEinvrarfTb7jn8CVYPH5XkHOgTHaXIQRQpQLXYbaZvHM9sqiNVxPoqwVOP
3sZI3gb3WMxSAF+55tN1pOp7ve5g8o2PVxNU0iUICUalt2i2iT8r/vMUs60veXhjt2qTCrJe9Jqe
fyNmqZrZ5ahasa3t19nTeDbwKyFXASuAtsqvSf4Rxnyi7MUHffW5bLHQSSlD84Kn8zJ+/tl1GMY6
CPd4N1Arh3tNbh6QWhWKBOPh9J2S8S9Lzo6ep+SV9TM51puy+Ka0e3iXUl8Pj4bQfQaU9DIBoEX1
HImQwqTEDhEntsBvxAqcblEEldCOpB7qRMhwpAxsGbh4Pz+qBe95bHA6TgauenJJ5TYEpW02ry7I
6yBRNKQVkKniPZVW9R8ro6n9T8Z82xDsF83Ha/wPyGADe5uUJ8s6sw+FrzLOwBdNRNdLbsvtqCCY
lk3bLnnIzmDppr5NJlJ87mhc0bYbLAKF8FeLitBTKmz9pO0upn4LilxckolC4gMWm9B6W5UYkx1H
+HLXs4aRm5y+77olj2W1z2a4En3Jelg79ofcoN7pcR2t8f48WlmQ5gs2rLumWKWAOQ1r1AUhSUrc
8jJi2kfQW27vPFRjIkZJO5+NJL/h41MYEkd726aJd2QQ5bUCbQz0mCjhrYa7pGvOnque8pQlT1sS
D+i+j+UpQEN4DewGsmB+eUHMvNDiqK5IQbJSsodGcu+vo04FbS8Cfl4QdHhTpZT52166DpxrHAYU
mJAOXJ/4XMXqDruwnieCq6dlGJbTbj25fr1ub8Xg7lPfdemsnZOqhp/0bDgrQ7IbyEmJvtqC4eXx
M0c7Pfz2o00kFzMGLBdRKGiQKA5OLlApBpT7OYW9CUJfRLHvf8OPx+6y/CyEWlKiHjg+HjV9bb0W
HisFFPPIfUyt1R7qLg6H3pxyWPl8g6lJ4arrx9yAqh1J99EDxggyswYFdA6rPwgT1hhm8s6CMcCC
Hw4OFzMSFSR3t8Elvavjs3rZxA6GNPDRihl2SeWiTfIEOGtdM2rwzCc10eWuuBZ8QN4BpWYgtGrU
TUL66xkpG9IwauNyj13fzwGnqYtWRpRwW/sf4nLG031rqnQcq0P6uzxrNtMNYVkeKpiyXsHlBGnn
mt6G8Qvu43ywxqfxp8g2kH36uVNJIHHmBxPlj1UD/f4FPFP/U/sW1BGloh02xZLEyRxjO+20379R
bEGo48XQeSGv047oMCwyQIdjKeHebm1DpasJp0fI1tc+CDDHrFsNIIlpypURBaQzXOlJI/fq/5y3
jU0SYqQRjuPW83Qnjo+yLJVwgvvAJFfONs7/iZvVvIGXU775uWbGh4ugC6cCtvOw21rF6jUNLrrY
uWfvK1xdTMFSUuRK1aP5D1McR+PMuKudZNumsYgP0a3YxievA5uK1okE/T9zUuLqkNrDWGNLzPrT
koIp8I3vc2DW7yWJALDLJiKb5r/njE8LpvFCQq7K8Y7o6B336wB6JXt0DvyWfJZrvCQ1mDpmD/Ut
OeMX3bvswQcNGQyYh3nijYgkg6WXpj1kjgpjE8FNQi5AQVDK4Q4Kz8f9UNQDTWt2Y67H37KgCKxL
G16IUOv02fazKG3UjSBI0rSTTl6N5BJZupBTP5fRS8iF6YBUUC37NQLJbVemu8JRLGQ/hCMnfZ7X
S7K0sjO3KK0pTnwqioNGTStg/MxGU5qk1RysSxIM/XKAEKPg0ebEYgNoL7ETIB/yIND3Pvpfzphk
wjHlEvbUof/4Ky5HtEet/BzbnpI8bz6DVKN16/+Aj978WhbEn3X3CgSZ4ncIhz/3TvsYUL0SAyeG
ADztPJlf8J+UYXcxNtN0v83cAtQNno6MWjDzCH624946hHWcJnKq07MhEMxLwm67thERrhIWR6Bd
aEGFsRT5tzSoyX6/NyolujVFrkRIUPtBXcepy887tAk77TDvK1qdxLlEd15QaWWT1fkIh73nOxXM
LCMUTcMx1Tzg08nCxx3fjqJPGXoEO7Tv0CqEsXOHALQfpVYr/k4VHTm2n1bcWZ1McFForV3f17tA
PTJca5e8LjSz+Q46Q5Se2SrM3IgiYEBDaU0iaoCh900x8IQgVJgmhDZcakn23fUrbwULyQrHHQ0J
sZa6flwg4XYnGIY7ea1daclaFLeq5j4qbIyLTTLez5OHAcY1I34JLAYgiEtXM4vjNyILk0aYtRjz
l3ec3DTHwnKYNviIggQZcUx4pjKdgKfW24pO+Z3tSEvzbI/6yXqZrB0UQYps7ejDDzU27wlLWKky
TkOO2ZPCahbckbbLOSttXqkIUVtr7ecUTD0arYxVfNyk/p9/KPJEf09HBMQTNirVvnBXF/6j8qk5
D7JxabRhfAUC6Cl8QpAGP7j3YoveSUW0mysRU1fmwwmUc9zDttQLHCHM0Hfhs7hPIohq+lHZyaWM
gM4NRS3Ia1khW88aow9gnYzYtRyCF1fZdrFVFsQwDyJ7YEty69tdmg7IPXJY2HNhEAP/0b8BPI/K
uFHRk35UUx/JRdEmbXyBrnIKctVqAL2DlnSrtFA9gJWb0MDJSwdldMHcPklQpINBJiuWssaO1zcs
HAs9Dn2fRQSgdWpcpX5gM0DlTvD1sQAk9lkvGf+rwIMAJxueCxaRx8ceSK9mrX74hGN+9K/CNh3v
+u3V4AtEc5cuo9U5OoMg2BbDek+tW+VFy5q7qZRbG7ngGlvc1C3hhm9mwCh2F38H+v3VbKxjLmnQ
gLACdvNx+DZgT6tu9G9sWjqpaQZ3U9hQ7ZspO0Y9IutwSuCsluR9fYtO5uwBA7dAsq9zc09wmbOj
my9/YnO1/ih0RGr1qFr+1VCIWbDKzuv8Nc92FbZRDaf6huMU5Jw0iYnFZLNVQDgCa2nqbI2sS7xg
zRxpL5KIQ8QcHPBvhqojQ03MnePMeDfe9s5/UrXigEVRaEmsQ7CljqfitI8GJnIi7cQYKesYav0a
Ptq6aY+2dQ51guWa5HTLzACYPILpnAZOe/djJQwMXKSmz1zj8UuVvF1UJsliAMF4gBGqnVJQzYG5
t2qwkzaUSPBblQy850uKmUuJTdZybdff6zkq4RVyi8jeC5YuEfXxqdaoTVdmqyMsNiwtWSGdvynu
TyAK9HuQw5mtwTuqoknIYzELOMB0EExh3r5jEOLHIS/paisPhIJdb81gnf/NjC7dohejzRCW0bpi
JnLUMCAE91/MVj5y/j+OQ5ZG7N/Qv6job4LKf2Knmc0P5+6NisECB1mbXzjmRI3Zs3Jn47FoGIEW
cSybx63NXV5KaD6HWI2njY+i6Tooi6M44xGseQ6EqXSVerU6fy3KnwJ4tiGLz2u0aQTM6pLdkMl1
2HlB4ZzFmvZAxeHHiBVBLyJSuPzBG1nQ/FAZ47YDKrqji9ZYe0ZtBbwJr0BEGSM6TBrkHjqVaxpc
in9bXJSmzhyVawo0+IUKci6n4nKkbxILn5PVvoMJ5e4IUTaD9E1P6XZ/MrTKMLmduaRIrcdosf6K
TV5x2gs2tkjPS7499UnkP8EkbNAON6/uZ7sBozyZggsBsJs10ktUZ6gfZtxwiDcyYVxidq9ZxsP6
LeSIB4wD3Y4wi8dq+uA3StjmRAbOHiKuwoLTBF+HuQdRKjF5N9JFecnOk+B6jeIR8pxTH0NHOX1/
KbuSLZLTcqEA7e+d4yDYok5qTexObxf17mfSaqb4RAEwq6ja7VKOuDpeaKATLqizX42ACdV9cwDS
pJ9DdExQAung81eh8oCu96pcB55zsI7HkPV1mCQ43dB1xyjiWP20wO5mvhINpZfiIk3mvNDe3KDL
GlJgsY/oJPXcH3PoovoETOk6yhiIIYVy6qtGBtDCYXmMO+/LInoUL4qU6c4Ki0lIpJg77VHT92lA
esR4AEfDFvOOzhMtsF5PkAiBP1oYpmWnY3YUlKILXIPYNJiAGjyrZS6WQhO/2SPmxCWRcLLNsTTo
youRNbl5uC5aRuHgy43mWcFl64dB7KtVjycFHmiSjzi8hYSHHxXAz9bAfYCChFTYvVvm8G7pic9S
tGgk3bLJofLzJw2hBXk8kOuXRC+MKjrLG3/UmmsNiHBIUJED/S7K4uDncHxN/fCSWZeJIaK6/8gQ
kxPhImhZRTUnh8bwWw0lyP4QoYtqn3DsHId3vU81bthWUX/S9tetCmdG39BXlHEIXp0Dh5Abr15c
4foRxDlj5oaDJ4Mf9bU7+3eX4i3EAiO1jzpVgCzRJ6xA8pVY1dCTDFv3hOZLs2z7yKaXNINFR60v
sbqumu7MkFCi5b7YPv74W+boCzjzWIEA5nbHB/I13h0IahGjacAuQ4yQbcXmmdYfF0Y6GGvrGGq0
t2IGCALEbOULA1JGc4PNApvq9uL2RXjPj6Bq1EPqzMnJaldBRSv94zABmM7E7M+AlNeDMt2s4Gi3
Aa22Ykmdzijif6RSjqJdYoOz4/T92gFI/+IejDI2TWK8GRn34NP1K7qV+X49iGU/YL4WRjx0bg6f
Gg1VMDbpzIFqkxzZg/CYN9umM31I9amqyicMTx2xYhzpdC/+hv+VBWlEXSPGv8QcAHQugQ9nwNSD
JABl3XsRCM4wadi+jsXflcx5D7hNc+TYOJG8oSlEFFuvrVLzYqPCYee7B1vOZ7FD9U5BNDOCc3wt
Wi4I3CWPDXiR8OwD9dfj9IbUop49g1EJYoT+Bur9crye97XYk1wJNbFtg/OqSIkl+SNSWLHbhs8t
rz5KIMw9QjsltetVGTkXl9GvURFBFYdNlet+OgsSSUpqU5iPJVauHrmxxMBbjSsQ+tAWKMJnl6ue
nqpmWngweHJeyGBDhpJt5KEfNG1YJnQ7a+qFCquwiVF2LyKlnYrdWF1aag+El+gcaOvF77kS33+U
dUpKIV4QMgWrIbWgfUisaMmBfWpwEV3mmCXzQ2QtfpIxo+qvCFIQZM9PkJTyg80tHQlwCQaar+wh
hpFTguizM0YmFbXTczGr5oCZrrDVkR394lOcuINKSXpaKsIhoNPykbAYiojO7n2YuTF4xynjGyp5
LShdH7VNEPmKQKywT0lYdJVZ4Zq5WyEnEmIsMb3UXy74VjTp1vzJRstkH78BUqTUJYsMJIeiqaIL
phNP0/2tA9HS1MiQcRI1Q/BAu3H3LfB9N7DgGONfQrMHS2E0aDNWu4u2rheBcLCQHiHfkt8wPamK
yqCMkOM6lCKRm2MS7rdreTm7nUxUo1+bxeZszOv2m2lG+turNkVFxF+P9abhqEdLff58K8/37+tH
6Nx8qGnpuipcOoQN/S4rsUgwrmFzAHXOk9v/eZxOBpNX71s/MbLp+N2Dg2FhfXQlVyr8JdYuIA3p
eB8M4cbpQFw0FcErmEbW0XIjd89vOg6PaE0ANTQiQ8R/fxMeZ61rurNr3A98pviE6QA6Sy/TtEjY
n5GAfBPVm6iu42G67BMxQPOHVXRzrGUtufL/EG1lsiyWSihqgVFEA9tj/kPHcytRxVTQibM69uMH
YRG5Tng13YeGMENeeLUVp2rGjmp0LxPKb0Kw2zAHR3BaMs2V4YtEkujJgAw2vPW31/rqck48iNKM
fpKI7ERUhP8JbsAWSnk1Zo+oGCkfHRzxg2bI7k2Hfaz7oE+v5cCleTCqCBQmQsgdT56Zxd5tq/bs
xFMR9JKhuP/Kg2D0zZgEJaxXf1wlR1dU6lABI+6TrvCK6/djSaiNi4ShX/s+jK+r9CoC0kzleFAJ
rvGjngAQucZgYkgEnng374zhabBlkr1LVby4f53vn36HUk/VldxzuRoTHh96fc4Jq/bye3CIv2Ww
+wecKuh1W+rNXa0nROHxY4M5V+LtsD6+P4acS5SgwMtwQmTSs57dSzAZ35ERFGr5BIMHh/k0OAb5
7uohmEb6CQG8YK3vMXfCiTDSVCHdhgo54P8e7IpZ5hK/8TJdCmnWd4B4LdJWER6nHOKBMTrmu7yG
dboCnYr0KM3nlfv98Ve17ORJkEG795AvtxjYSikVE/K8jSJXuBSzC0Yu8krtYdbsZJir1K+ljuFC
cyK4J62GEYMWz5nel4SNKVFhzNBLvtd9AgmRmgGRBUTaOkuC/w8+bMMz4GZ8XooL8e/Gq7F2fbe6
tiJDGKTVB5Ssu+igxPr8eYdbIHmq58Y339bG5jcWCAuj4ZXUFCqQbE35LMZ5KBJoMxn1gy016RQy
udYbJ2tI7sUchbffaEfjYmOCs8Zltp0OmbfZDwHO++Bu5eG6aQierVnmWx56Myln9ge5VGsDlJMy
s0/zBItr48BGmYmNypXq4dgTX6r7eF6dnHXtdBZYQuUjirAZa/VpoKKOeSdrPVzwjUeBoq0XIoIv
z0BFGKDacVAGv1W8NTB2A+yJC/8FlCopZey/IsyTw1zWPEDbWREO0gmRMhUXtgWuPdmlofNeZimP
eDvCjjScAUA+uR/TppzzWCsQM8WTRVJHBxYENEjxg2Q7jjNonI+ddV+FUbXdcO678hhnOeZYWfto
vzoWdtJd473nR7cslc3pMSGlYUc78YXs3PNDccTS8VUzqNt7vhArPQ19bxYjVrA79EaJOTYKUsrK
XN87u9f3wAy0vtrZK4BLrrNI0iRFSPKvh8fNPQeCsbOcDX5bT1txUoP+tItFJDLUeGzHtLFCW0b/
nOLhMDMIFtM+oAIvwRjCXTOlL/co7OxEJ2NQFF2Xisx3a4eY0UyGDrJIksTRJv3A44E4QdFa3qX+
7VcEYtasDB1QWA/QFnNtRh4IcLkxUOdLG7gSvGYexoDEGfbLPQHYsXQxNzLdGGpcoUs4h+CktN0b
1XwtQvlT+Sk/ohSCHsXQ61BQPxKtdGEwxILT7+WjhicgvnIjhsPIWpREjXGrHVcYbrGvwJzZ0mpA
F7L/BmmiGfrttHNGXry0vU961ju/U84muezu4bcRfQT8oK6cPMRQqbMiDKzZecllaZS7n9v1lhrY
FdI5PHovb1fvypww9BzaMpYapEzezUM5iHFAfFJbK8XLI9T6F7wST2woRwAI46wNAtP1ZrrcnJG9
2En3y15Sv6HfTY6G/oUDAfEgaqeAaeKaiK4V5wLWwERn+IYN6n4M1AGeJrDl1BWpcMDE1tt0PoNk
CSGhR8BtG2xUK9f9UEhAnQ0twciuz8oidDTBRb6kOR6sBYXxbfV8V8NTAd9kWca8ubFPiOhD6Ro+
l4zIG2aHcXznIfAZ486NqBOG9izKqLow1VigBgKLMmgw45I6wnOAgXDFjbtiVFxQMCCSYwJlQVtI
lMeTVX2oRHIFYqHOa4S6YvYo6ow/SPj68k2uWLz/xel8sdGoeGAF2gjlikVhafq9qo75SN1582/F
fBC++IpCEOVZK9CVL0ausrWGid4dPzyzqYOCxvRUQI52Wm6a+3c4tFl0xM41/mhjExIX086WplPa
Af8UCRw/8sU0rdTLyM/6rTBCrJhu1EpwqvCv85uDQnYBP1Nj0RpCGHSzp7GlJWdi/pUh1TfeGt9A
nrpvYCxO7t4WpGP8Rwp7JJTf+GOjORzZokOTOUcaiz67aKSDYYeZr0mK//9TM/+/FPvXdY44MfS/
H9FHm1f9sTzxGZAwxpEmnqE+UGngO1NA2rW0aHexp2qe7kSpAnskfyezNeWAx6cKzot5EvInTNTS
wRK+Sy5Bs0MLdwKVdCaud91mwFhAzfNWoShpKTY5GglsvQtgOJ/hOAS4GGJGqj7yekEjhtxhcN2w
TFuiM/LUf2tPA1BeoTXzRUudUq5NF2ni8j1Vu6QlYzUCp7NQjJ555S1t0kHPI5+As4OMdmVJRV88
KJce3eTJhE3TYV0v/gGPjkLroakQqZY9hLbrvUBT46bLHonuv8FcWEB4/qP9u0om+v6yFlIIorsq
CMm3MRfVwIvGOYjdqmFQOx7i14kR7iOEh26lbjeCn1wzZ4GD7TvCdG0mwnSGtXNKLyqzuzpMZPc0
yRDdoKqhUEBYW79oh8CQd1fZO0op4Xo8WyvfnH1hMh5DI68QxQiAzCRRQKRyKRDri39bswZaeV/5
2W4yeBS+INMQZb3otWMQr+tvHo0bDfyZPYGTFTwwpBMjsM4bwWemXD+6RMeu1tdWHQKppCXKwyWc
A3RvyY5DhQR8stWY9odZuUrW5r68IhIRsyajOxzX7ZnnFRz/AUc7rZunjg8bTwD+pziL1fvRUaMc
yO6IU4cl9tIkJz56oLpaA7YHGJwPK1b0AOcHZHtO9nZ7bQG5zNvwGBrvC25X8Cgr4GJH0EkFfqof
ymtSeuLp38DLyZQwVUlcWClJfT1k7OzFiLUVdzxbuVD+n6NAlcddrrExQuq9NKlpkL7wApXAIiph
C0ahHjSOjvgmPpZNaPERRFzSmsmN9Ca6LZPwKOUca6TYbagDVxGfuxUk0cM8QhoGqq/QjsRBiXxX
nTpabNz2qcO2ENlR2/I6wiXK+eoo1RBfTuVtYwJNLfJfknz8rucgpcWi9+KDaFwjWSl5Imxomnyr
1+DF0qtz7HbhaZ4rG9IpdfBL9N7A4J4sQdbK20BwcCdcMrNbG57bxDMZ5eMdNuKkVt/jhcdgQBNZ
xbyMOmWKKQY+CXyCjJmt/G8XzJ4ALEzg5LnGT0Eb2lIN/3NgkrxpExBy7INDfFxpyj9x/4e3QyJ1
0ixnQk4IUxM1YDrYIn/DykYA5/sXbfAHOwU8U5qaBUmbhUPqvULNc131DDsMos9Sk+WB4Y/AtCpE
67kG5v3TIn4a9UnpSCYTVwcKQAJTj6BUIV4QAbgwu5cVEI/tBMYiske6Fik4WHODbFGVS5DS1Mi+
4P3VRckAPgxGeC+ehv4LO1yskUpwLVvyOLwmgAyXdUXyADVZsEO9kecPf7V5T5c/Ler+6Tfm1Po9
T5w7WmkKLp3w9+vII6zF5KPgmBGy7aDJ3AMd1VIcZJSXZcBnTxL08X0WLVsL7u79ft2XtT/H2W9w
1q3zMcIn1RQvDf5e1lO792vCYixqdCHFZz+ZtWgdf+J9UM/C1OQrghYhHr6dW7loE8R7/PR9BAaA
7zsGkTHBPsr7fde7T+lxB+IehU5warMuKX2xDo3ALczT2MNf4+sLsVjqbWQnK8RP2JnY89F40vND
zg/Qtv1qFb/z/Vg9h6tVJCHmsVtGWVnWPMomrm+PtiUiYFc2D3Iqzv39GTGA6foY4rd1o9wclulQ
xQtACHoCu8YMvCMFhuQtxYqDC/fUYs8GiFt5eQgSezKtvmSeWOmBm4EhQftMRpxU4f/RPRSW6jip
WPSvm0u2MMsYejnZJM3qFgoY8h2PPO7DX7NuT0AhxknWGKnxgjwY9ASIjLggEPM7EmsU5eP1fEkA
C9co6QzA578D1JmWVpYDZG9h/2IsJVjOzOjgL+wwKyhHJ9fop5fgLc8HaW1A7HaIEwzT/UgFXCOf
zPRUnndZAjWwRHm+b2Pl4UvKfjLUyqSTiqcxMTNKrcObvrVS9imxHgA/wX8Q2Lk7Gok09qFT+cy2
h2oKKjmd572dGMOh/M//mVqhkCiR4X83KqJnw4iTBn6ly1fUfEbjyRdjQ6x4rwtLuXmHnjhejLsw
TwtLURL4+QKpAm9H0o9odbV7t2lvJ3uUqzYiWO+8SXBWTjMXv9QQUPex/kuIJADUTdm1EL3jRs32
QJnoktCx+sRBFKZWKE0rC0pu+25Ehak/ioUot7HOdXuTVEefbS8AdWIdQYaEgnGhQNrMA3R3D2EX
y8zfUkujul4ivEH9sQbj76afMY3sLh71tbYWfkm0Q5R4HnWmdMyMBFvhhciN3PVW98nuf0uJk5Y9
1v3MO0+Tr6ZYYysVPq/hGXCzmppiN/WWlYPga8s59uhC6TgMpbjD6MXRJHOaiFa1xhAuzXPGl4xn
2TdAWamt6ILK8u/VdIL9bPAQCBlExSChkbeIPAFE6ZXegsXkAPSLYwbRsoCl6KSsC2AgYz3HjArd
bAYLJvz07d6O1AMthspcpUemE4kf04PQ+3ZFLnmq30ZaoEPWMq/zFQtf8a4LN9LMZb+7IXZbFTd3
Maj3NOCfdlIeTcVvhhIcLFBgUzzCbPMqNdlu1qeHqfP5gBczwfVrzMP7C9pZh5Nep2BMib3FmvfG
xWNUh3viyyhawX3WImdT3iMzgMJ7OsCCpaWfUVqMzjbLEIMGDXWoae8kJc/XLzP2Gf6sL+2JLyh8
/cXSqktgH6oML7JYxl7u520Zok2N181/ExpAM7YBvDi2/gi4P19mG/g/YGkmK6VoaYeuvK6ifj6k
fsmrqygGOWe2wnnnpIM04hxWPn5g2g/iHdqFIVMuFdD67eSAZnjSeeSy2etc7W/q9pFiw0DBG4/7
Xb9UPujCzySwPZrdcmzJAJKkrCXDK49JtWrj8WvBObOf74L7ch1ninR++RvbvdGSOB4Xc9CmVMmX
a24wWKVU4sM6odA++a3gs9ZLUNVep/GBAJ7aWkx67/dgo5ue3RQ3V5bOVYpfYQBbyuGb1cJ9CM+C
WArWQn3OUYlKGczAN+HSqfSOw6qvHhfHbZ3RAU4U+NG1vDUszWdYadvPg4LapYuu2h4LMoL1/1r8
5niHfffzkfzEqBPOjgQGcbAU4kqmrC4iOre9eeidm5pyPv0LLDbqGh+ApvRdHBSQRsp3dw8hvcFP
gs+oPphzeihdCUov6bdOIdjY1hczODDClkFjAzEad8D86m1oV3wKkkEsqVT7x1sMdyYcqLtxv6w/
z6jDP/uR7FsnCJBIzI1D9u+m1/t/t+amDLcamgW4Sdo4Zc5urX6iTCM6saDrBwNSjDw6opNr7QOY
v5ldWAqNYC5ObMFHfK7OofFdR0PPUHus4plVAdSlwsmHqkM5rB+YM3UbG+X2fVwnrUHYxkhnaZYx
YtBTcdzX22pt7wYmesx5GNRHu6nhqtwyBVqM8YC2l85MTv6in15G/Y2ipcoXyKEXmCIFJcxUZ4S9
2mNWGHAzoxeR2DSbuBAgElonoo0nCdBCJ7YHQVErwmhhqp6CMf+/Y8hfZypPy0xs/nOo7AYBel8H
y5hbEBY46jRrnA9EXgFfG/0eC0tgTtl/zSduePWBORJvrxS4lXYB8ysuBQLp3hhpmYYiq4ThpwGz
OFzX4rUKPjxwZornv7aNkKyZ3CwDQHkjH+37lrzrCxuR0fxr5nqvRzf9KFw18jGKfiBJo8IeQAwi
ngk4jOeY8MJFJXFpRJ3XsluhGa/SWltzwkAEI9yVaaVg/fgsf7TBlPmQcMip8D/vt2+SU34dIqLn
qMXLCV/7aO9nR3XuJTqS74eXQeYXldwL0YLdkEFivF0J+3LtvO9EH9aBwohREpUhg+vGLIdClqyY
DG4z+OFcyaWfLfKO9V7r9/Da6ExVOAYpoVyDTf6MKRkpZiyANu+eKHUuZ0tg82jbtl4ase15T04V
7IGb1EQcws4GyMrTwu4fMoIXpYG6KwfVangvRJ48m5u8nMAXxymqv3y/O6iT2FEsc5zG7Uo1aLJM
9G1GMX8lxTyPER87bfPa9kkGiVZT9PVY9BX/yIeSzX3Sxpx0ojPbZvHar3aywDRIkcjVtxKOwJZo
mqtt03UUuA0cjcBRos28DtX1gV8EhJuup0OjvKrD/vKrvaeo7lJP2vclP5qqeUhaoBadByljyH08
ux6txBQHF1MvmggNFfR7hfVqt2sCLMA3jGyLR9qrsP7K1wUwdJofstvm9d0f8bn8VK0mb+hW7Bpk
rLNxFeLwx2v16lHRFVD4GsZlUodr1n6ssuqSzOTywOwU8MWh6EeAEJSc+hrOtC87tmV98vQoTKTO
3VOXsgpanvDGZPZomXsEeQ9paMSkWsD2sGzbRq58Gkyd1SiUOzm7KTRPeIdk2hu+OgV8vTHm/xMe
op16ozgreCFe6DMCEjIL7wKhP9dfN56/TIGw6JUT4mkWvHr4eEZEicyKd7xDNusFRimrlPTu2xIt
Shb7PzIXD0zt+YYEPRk9DFDYsv2XsD5nf9SY7IoOPPFWER1ghRry4zqyktc3cu/ou7e7QKrlK6c9
JxW7OLCV/gfYLetaqRPjxmTThtQkikYSOxGK7AFeiP+cuuSKeRec9nKlKgGssz53A37fJc7pZ8pv
a3CiZOmFkXEOpTqFORyogEStuXutLiAiESEPFOdxiSBiRopXVxBnQl9Via4e2D0r6ixEqvPnY6uD
o7anog8oinP4P/LJIor5X69dnoocR4ah2tgfjDVGWgSOVgUOfMnO6fBLrscxu5aVXnPqsUO2Q29t
5rWLukU6cus0Ype3wURn2ZtOLc5MhixFnlVyh8gqrbABkj8ab3/GddhH/Yi4ke9i3t2/jtkGsNiU
rBzR/hbGxe1mj4bPKvGAkOHl8FFX9+vFBADNzqzW0AuDyokrRMw2gM0apJwqEdWxQACCOUSfcGhv
urtskIJl7U2EA/9ovDqnPQ4S37Q3GrsVihcAHRo8iVrmKFj30ajMhHQSwd88eBP5fsxv5CJbMQud
P71Vc7TCHVdvjd8vO32pjjc3y8OyHsUkmPwEAzJHqWcd35qtvOgAIFV8pg4EVUyuOr459crVw9vz
Tutx482Bgev27QHyneorJmyXMn8vDTnBmZgK6TMY2DRlRnAMxMKRMOrjDM20MsFbw+C59nkR5OxZ
AgGGWuJgc+FHPhNxhyVg0PPcMqJc6qQ49K+Ady9pwPQlCw635AztXO/Tm4JQB2pzZ+7zg6PrVatn
y/LUOtxRYejWlDXA5sw34X3YJIvOUvTjPhU5MqWDMDpGCcX/EcE4ohZ4kQA0iPhfvBcGmAfRGsD9
d7UYTxWjw8nS96sdTJHrWqAurqX631xiLABvaRh2vJdV/CGbhjtRbVWyB9BhOcqrXbOATRVtHJQQ
jsBDbZL+NNuBeTI7iQKEExRQVNbY25I7PucfI0ruCWJ035rTrHGRbrFAh72OeDtI1qHGCqy3oc4q
tGn5XPd6BuNz/AYw74wwgIuOIyjE1yC9jBDdV0BJpzbr27iwuFq8IHl4faMI95PffER0akTShqYJ
4TpaZEXvTQTsaTArM8iSKVDwXwOetxfEkjk9oRPXqv+KdB5ol5w4jlhiQg3R9CuTcv9mgFv+Kgoc
Zd7do50hNujjHyBhrLJ6niSIEuw+SI3/GMeCOvjUmpan8JdJdicyJIog7sE6qImvVFPVPa9rMZ4v
is4Yoj+AKKgBAVy6iHz7e7Z1oeTXg/0fIKoxBOio9CgXomV9ysIZ+IEhC2pRQPeRmI9mmBPp4gR6
2S8ewZQSZlKGnZgzDz8qcp68RtgEintPV4eBu5OZaN1g6P95oL8zw0xqGlYsqPwToR9rUoSUWWsv
QB54UeGodIWa+g9uk0qpyva1ST7swvYNYEK5kEevQHE49W5rKaCBLuIfacCPjMgJgWxvCdRfR+BU
ERR8JOaA2q5bzKmixYEtatOgk6vdPf/sc2751m8Cbr//ad02ZAip3D1tESCeY1MTJ/oN2Iv/S/11
9pwkHZXgdHb/3WkjdMgcBVgvs6LXSVdszqRDhyN07EkWBMdU1fs5ADmMbrz/sLoFiand1oChSxVH
ldrrUeHQZAdmwNICFVXNnc8WNefsUVrFSIVp69S1NBLf0I1XW0Bad8mfUVXpY+5dwv9HZOWh86du
ZnGrTUnjIYeNyPYldNaPp/+r9VyhRyrNeiulwMxWu/FYa8Cm1l4VQek9QMT9swwAHT1mqZh0Z8ji
e4kuJlRubyWJyftMg3nSUaQTDSvmXHvh5dmjq3wWhu6Yj6H83kzU6+akPDRq1ZsbkIP4sx7axz5H
Eq6V/qm72iVPOTvOH+dX00wPLnTqMf3CB6GNvFf1sUvibhoiokLiHLbLYKCGwv7ow1+Zhzm4Y1ZT
qdugn167e+OYbblprFSSMLRAunQal8MggAox0NhJHyrFQwuvWHZJ9aZI8OoKPudI3ozT75k4y3rb
EnT3f886F1+hfBJjq1S8PoO8/ThBoZ3JZQ4US2MjbdXnn1Q5ai+ZhmMNhaB9yxVHs7hufgtwZZ+P
DHmIK/036ulzmt6WgjAjkv4eAy8gFYnpbQ+ZFSTEO0p4jB6fF14JhUz5fXvqeKtRUQHtp/zAm2oe
/l6nKzehmyyqkRaPnoYkxwODj8ysLiLDVy0HOJ5vDqJMHvAMhoaaHy6G6FJA5zLZZ9SpUtvUCR90
VdkOznzFA6K6Ysr1Pqc7WT92QX/+JBLXtPp6zjISCVnbVw/ziglLBRDYjyfK68/elyj11HvGJHVd
PVBgT5KIx4fy+NoU0zbKVYcpkoNZtSYfq9txEul+xT0cY6y9gA8FrCkVmeRHBT7lvjEdm5op17kS
pxgc2vTWftj9ZY9fv7oOSvhPu6nZneLCVMPeP8h9TsjLoMcA0ophDnKU8zpDDGIAisYUQo+x5qJs
s5kxlzfltJcQC6m+nkqUnA7sTmt8Y1j6j6cs6lBJxMj8UZsWwKaknd530LsqUl2o85Kyc9YfP7vW
pjd9Ujn4Fb1/8nC/BCj3Vtx+Wu+PaKYtrY/2+nKfSl+9Mz0Np8R2xqxoDwci9KSXN4kdxh0jHhOJ
Z92ZcYPOmiJWrE8sy5kbEUBwCmFINnFxXEWg4jbky54esOT/uDhRHC5SzrRdfGPI5asYDUo609rA
wZ9Um3iS5ZvH+TWPHeGjFamdD5HtcFxgzz6tk0BCjdwr3j0I35KIJkPmk11h8X+OMvFEXlXLiHNS
Ltzum42+UHCuKzKi4+k4Iki4qPejnqX4HAbClbFNk1EXed03F4hU6bBYq20vcbqiAsyj5ggItBfN
3fPz9yCTbF2322QRlVoQTmHbECVsMrQH/QWsu2GXX66BjFqPDquVG7iX06j8CYx4k8QWirWDpC03
hxZnbK5w/RfQXdoSl3NLQdLE8Jyd+t4zFCfn8g48B9wL0jXKwhiXPqsvL0sg3/YkiWQFeutK8oTH
lTE6cu8J+NUxWf3SZ1KyKtQ2JltEv1z649IkRxBQzci9KP8G4qMM8bkP6q912uiHPY5L9QVXY/Ok
9xcp6q6cgLekDqDe/qtuKeFYW0PHH1Z9HrmtXECZ0q3//ZNxOJqzccmm/mFlrRU0Ly2i+kccItYm
NyzptrMCauEIVhg7V9qZ+0cgh/d6lFi9MQ9jiQzABuBF505HZSCeCqwE3NBxufdvK7vCcHZK9yzV
iyVnnnQHO0RZl0qf/RrwNoab0UinYrjTaSk8AdZ3KqTtwtLPSSOHqWNEhngwN0GVC8zDAONSwaXG
RKJbAV9A8s9yhzjHZvUSm2aM1vx8LfI+JWkEVVk6RzD/TKWJcfpQ2C2xHdkqePWbIGqPtkOfDVSt
5CDbNuwA7qTCkqOYRPicI4dyY5/QgSTn2UE0L/jfteLRpuKIcPvWIqy18rFXZOs6DLMt5p8NNpq1
fy5Jv3W8vDMFc48ILX7ZAVJj6EH2Gq/SCDDKjBWu8Y9buuBCQDLwNxa02lQtBoUeUNdTQW2j1VK2
wFOlNZagKWX2n5CJi5ImxDPjo5Ql6vE18sCoc0x/Ak1+vKOYJgqmm7p07QI1IdYfpMloLuwTkWDl
LUO3naQpwH48vbrSpjrPXGEfDF57h8IxIzPLQbEc9i3GsNpmvANK/PEDg+ukcRnMMMpxitbZ3SlH
xPs385eJo64mzehu2+fyPLjUot8mcLONGMpjFKvPxRCserXeH+Ple+in7Pbp27lwe2YHZYl1UuAV
LNSB4UpGFRD8Q25PPDna12gsrYzlKygC7nw/bCwvjq05huv2jRtwSyOnc/HioMUDUKGV1Q7ghugj
rI88refLWEIozwO8dilE3jCYLWzJrVm8BDu0IBHyN+aQ9GWiwI8neysPFyidN3Uiozf73LqqQulu
b8pvetUqT8Tg32WWdxYhkZxusXQeT938oIkgI+KL1SLjfHuKqt/4e2s/sO9X6Kw6KlmeavoHL9r/
mbUyEw6rMvRZ20K+ttK8Xkz8BzlOhlsG6hHAb4Cvpk1KI/xmyxu57DZ9DWJbF0c++OZM19D07faf
zIXgWj2Mh0fB0irQAdTviUHxJ5YzpmccTJn8gH9tJliH+mfcyf9QqjmM9cDOi90CrlvsgvbU2O+S
9eT7pglK3VTuuf+70saTYDkvQaiReWE1X+qT2WHAjTZeozZ4oQSMqxcd1QdDSZiF3MMbBgKhQzJZ
S67h2kODID6vu9gZg57K2ohb1RSFLhf6rlLYdOV636ltOigexrReGNa4sOBlLbonYwdSkoV7bCmc
EEIyoAdqXwOZKWKrsCtqtBvXy5lH1AM9UyhcldY0Ignzryhwx2YNjGS57Gan9uF4rew+GpU6nVSB
ZO7nYv55KfbFmltjfHmmG2N3B/rWpCdAq+eRQabmBR9IZyI7ulZgrGRCyGrmRclC2UyHgfyaG74W
J0xkcZJji3E2MJhSCHKX2o5dF6RyB7Hu85IB8niOyxq2t0mbmZ9a645NdK4hBW5bYk8WvdbhdcJN
i7IgOG1lm1XqOByASqS5YyGyLuWE8cH/3dNN7JQ/idTerrIJHxZ7ujGs8LRXtH65Yh/FJ3DDionQ
ngxeCwG5RATH/WpgnXRMRbcmiWJK3oUb8Z93w1ieto5tY+Z/D5bUN1mr1+P+BN6vFp3JELrng810
bj1BJ9DP9yBr2ShKv9L20rb7hsWBgJjALZl50ouNDzwE8UvNs+sEUprKDwBNNE920V4fMh52DBIu
m521pmpF8LZh8+t8fDnMyngrxbq0zqbuG9K/lCJ3TtaCcX52GeKzPpBxVF2N+oe9M0FAvlRBimeh
3OROqaJgZpUSlrLpWuY+JO29ZXShV3lTSxN00TFVY3MMBpiWeseboaclbhFP7Dxv6jFnKkRwZNcf
H5ANTO40TrVDo7u1bJ/mUm1BYIlcOlDNQ+SHwJpQQaudj/SfOA5qYUhvo/gLZ3FhXSj0R7HT9h4R
rvJkwiMcbC15GXAqvb1vryTJ4wp1SD9W3gPMNWdToOVk0ibN+dd01VdTsV3BqFv6UkHNZ6QFYdqq
oYt0+vsAFLJe3POVxb9O+oA5F0H+zmmUaPBit4T+ELAaLkhDErZdoGQMdNXEWrpeiKG22NXMS4BU
C94TkmxPTsYRKZbrc49ukN9ikrKe0cM2JV58OIQHtJiVJY63rcFB9RhdPDzCLCEEao8YHPfWV1/D
BetF8WgKEzR9C1h4HaU5ULLchbXZcY+TbYBHAbzlQHDJ7c8zuTKBz/VHg/IHUPcS0au2o3/J+Q2Y
yjvNejuh43o3U+KNlltBUkVExd2YD1roIymmRcmsA242uJ8fNOrbxHUv3V2zOxHSgY3LaxyhRtV8
gy7Xe8mGXUL+d1NZL6lhpvHhbL1yOZjQCmnnymwpuNEfNT3KJhc13uwWmrbIL9GHJxjmycb9trtc
l52Xm8Sk+q59CPvseX5jG82bTad24e5/b6CpOb5iDvVBMOGgZU5ov0aN3oh7Ybi3GC2SwQjEtdHV
zqmRaBKwI/XEG1YJ9uoyxmftqUXCLNY6KacOP3CPReEFj4sh0JzGlgM/Pz6QGgJpK+Xr4Sh7ibKg
Mz68Uukim1NGVkig/NjFGn9nJPImz65aqXppbzIEcSqulziAhpO/21pXn7pOmpsfGoqDbuMy3bPL
QyWbnBHuAXYytBT/5t+wuaxzxA0eVjRLKfeGPB+wIh3iO3J4lQp0XrQy3n+QR0rtJEA/qWDfRt4K
gC6a0NxA+cq0ypE0KghCJirFcijf2j6FRizv+M+Rven/Jpl6634wiI0vg7zffPsTfy0whHEo8hOn
7pW3erNap51q1rlHz1t1AuRC9EjMZT4V5PctFTRiqkFfMBz/FYlRjwTKL7IWPtrmbxPg7zlfEH6V
dCeA/hXwcSDFECBYrm6wbFGlN0mtCtc5jhU1uaG3HlucLdvSELkhg/6SssAeKVRBejBzUWNVdWiY
mLADSYBw3SauBAfM3Erq9P1iUPvgrs8BUoZj1WT4fQ685hIgVyPRQmDD/ffpHYX1bBe49fihQLHW
3qcaKQd+ed7pzeVcmww8Wg/fahszrfW/DI/uVAyxOktfEiEyO5jB7B9cAKKAlcDxC1xG7KNjKITV
SwfRIDGKVi85bwNx6fiEkCFHCaIu+cyc+P3gVQpHHjToFDigrNFgCIt9Pd9bkYt5kbY0MjVtNkcw
WvHxv+KQdC/N2mu5l0FIIuxN6JtoG/EDEYQPCzXzLjGQPr4Uf5tBePmIvj0vD9rRq//FNMzRlCdN
ScB6qaJ0qyMTnX7OkGK7c+53KOmfUK+gYaEF0ywfoI/r9J8Re2C7jQ90owuNTHoLvuXRcMncsCtq
mjBYoxfJNL0dOm6gayx8Cqfcsah4bBxJLrFXzUXUyTJm/WK/6SN28QhZQgjANLHidTooj0uGvUaV
n0iT823jWfCOFph0muS8gENkTwVsxkd3r0ac/1hEPPoKinpMKs7sS8TixNZRCOeHPsaOefdOGQuN
QyVkpsAT+W6xyqJ6gv8eOVy/nOincbmXWP1qsh9ZnalDWyOmuWp2E96EjRtd5TyIlBQdlorJMN3Q
c7R2BY46jlzofBS9NL62J/8hmv1908WSfg8foZukwH9jru4lBtZb7sOqPb8LHbdDD4xFkIu8sDyI
g99zKBhcOz+U1fEMYBWvN7PCspzoBaBTFwY6G3cdRMOWJcF1aHuNN7TGgRthdPNaW3YjGqChozkY
EfQLgcFsV/O4kFpTFKkQEghWdsre1dyrGLHca7HWex2Gf6JVmCq5VA2lwIJn3kciXaIAg5K8wSJO
VTXoCJm6I4crNTObNZVVMm/Hl3v7SmWM7se+nBQG6SDmtRXhKxHXRtG0JbuJg5B9Y5jkPPyCTOjk
QnUC6SiUYNQSH69p95hMzWTF2D/XXMSkcm99u8HD6fbkHO1QfOoc7lCGepgsjVanNGoT6l6l8F0i
dA6HhmUhBKeBwcBDhju/0aQl5Q6arJfUTtUJems/QEm0A3HcC/flmKuEOWppj/OUK6Bhg1sFU2kp
AMj7uDSxNeFIjMNnhIEP9TniUkS0fKQor7yOo1grZ51fOVi7WsPuVc/XCAo/tjEM/+62H6DmOAVp
FDNTEOXb8HrWc8xd1+mI25bpSjmXf3YHHtyeBEqRue0agUzcPNfpX4u8Ii7nWCd3TfSU0OPB8jec
gTnqXWW2B1xIG8IRBvNW6n3rDcWG0Ilm4wlkgdlZ8f45AnPh+lGQA/JDtz31du91H0151/iaGhvW
NDYjagTH3zUjiO0pmrOguBsOWcTJZiLT5d0UxW71khhUSyTSkNqdwO15ZQ/6mIXyLCGFwGhMsBuB
9jwPEH49QWZXW5fZUq3Fvbtckv4v5ip/Jajk5j/f/m1ebJwRXSuU0Cc70PbXbs1HThdyrjWU0tCr
9pxM5SJLbxsWTqa+r1OzEAgEkCBZgWIM6DvDAyEpmwM//XCfCRWFQjdnyy5XWRz1SzMGS+S8ktjY
rh6U6naVmGNucANloD/XvU+TsfrJxwlj8N5ieNz7lidt/ZEQ9Rx2BJkbmiGFJ2W885oQFg0YuXYH
Ui9HHFpZ3fPzp3crQ5ig/QE+nVTaG6oIsf9CFtF6IXszwipOc9VQeZ07P4eU7t34/nU/WT5vyUI3
OhpndfJEprUT1ZJobVOtPsv7lZfBIghcMp+wcOw8kp7kDhMN4O1zKLQjN+R23VOhnVpZOIwXoeyD
gDM40InRAp7e8jeArvluw3/SdwW7iI8IGZGY3IyTk1yQsw5mtmKkeYwmTVgFYwL9MCYnukODuEgO
gIKqb73yam1hWjUvlDqwriIE5m7znMLcqSN6Mjzk0RWcgih3meHS8pgliamRiwwGGbULQzR2REro
Lm4ZtzYCrOPrNO/M+1sn3K8qyLpcTdkGUULQibZGVwpMxglVA1VzwXfFeDl/f0fOjQb8XIkLAwdK
DR0lMRKh7yj6Ph2e6luNsOFDoOSQKrayBih1+g1oxTd1em1xX1EDMHWVD7uEfOS3Oe4BzaRYuL4k
419JaHO5zh1fUhBwrDBIJ0FKZRUvCA5kAnyvimleOVw5lLkusH1BTrKbKjiCIgYmXBO0QnzSx63M
DqrNV1I7n7dKvTK5vxJzV2RZ97wmXFUl23+Gwt9YFuNC5WXdz/e6qPumY8nx0hDpiozGXY+5Pu0D
1JPPgRGbehWbPLDEImGyiYB7K7KjJBafZ8J2/YcJc5HvCEkFqa7pLH8wPpeEDiUw+GpiEMo3NKhN
zh9qbjEm6tuMgaEgw4IIGdMe8HMN0FZCjS8pMGaeWfYM++wzJLSBVThg748YJs2/7ZvD3dFoerIs
5PuBn2XPB5sKhT7+RXxPeZmY+KHF4Wx6l895KIwZP1TMViYBxbEBZs2lYb5gfD2qWFum5017TYIL
gZUM3ylRePptuWU9BPeCKaqJAi+3fn7ZNPtJSiCN0Gt2aLQphhcus6a/p9+JD/oI6o50BiGReArw
bXm+BZ6ohBAwpmvS5p6uC/0rSJuZV9cW/r1fWTq8Vyy7q+bxdKK3efBJqxnefMn4H2AWjExprWtT
4kPxn/Ce/Vj3DE0RbH1xMW9FYvWRvzQUYx94PJO5CCrN0gb3pjexnH6WBMilgy4DgO4pG5trCLN0
X+ksLWplSZr/k0lJeUHTmNZJh1+AvlLeqG+0mwAgCrg1gvmxGHmmfo7KjhaFCPy2ymLcyKnrDAja
qIM9yFBbtGdC5GJpsulQXGe9U2zggQs4P/sHx2c60MA6LSsHYqTnuVQ1U14B5QNiw5CwCUyhVFT0
vHZJdGRsercPTjs/DhXeZSvfUdXVn/oLNGH5ZJNmyJ2HzgnGP8ABbKx3C63Rfm49LTISO99PY4/j
aY//mCkR8p3nUMdQ34b9CAk19r/XqVHPjy4k5Uwlsu9NVy+BsvN2ESrayhFAuAaOr8fM6wnVyArz
SK5GuxOZix5uhQ+3x6XAUljptXSy0NjyDarUgzJxxB/4oQNQjYmcTN9oKKphV3gpCPzfCNezXVcL
l4rDfnhjTCxkmnb58pqgM8LwSgkvUNRp58JLfQL1QRJOe1qMw+FEN2ldhPXWoAVloPORWNPTq5jH
m9UUIbRQDC2oWhAXf+B0wkFVStAwfWgycN7IVO6TghAf6HmIFDzTxUSez4GrjGT5HhIXWzD388Xe
6i27r6h1hZWjq8g6xKZ6tBnKkLLl07dR0S/FUv+qh2w4mh5/e/z7Esl4n1K/WKC60IVNh6VciP35
N1/vvsB/4fdU+6cZ9o8OAbF/YFnKUkqZADEib/ZxKeFA01hEbvvVurjt/8Qiaa8TL6/XaEbGQArB
LeGz2CSVl+Crvey+TUx/8tDQ30OnvZ75OdjALn/vHEpikbtE/qJimi/yNEYJYuGw78tcZZIECVGg
koHJY8Lgy8O8MkJLxUwWntJsHI63vYbSi00qNgQftaHV+P0Gav7W0Zzjg/9Zw09kPEZT40mzdjgr
fn3Wfchph5irXiW7pVTq7hSrezSXRko19hcJTfkdCbenlKK5BzS3WYziwtaAK92IljM3wy1YMFV5
O/fetRJSBJsNbQM/sfR36DGeuQ5dbQ39CoVZA7sJ3xDoRK/JJHuoEm7/NGLyXMF7Jo8pXQq3lUsa
Onqz0SdS56WAjHZN+pfO11j9owTL7FamTZCi20gO/RsGskSZjotm4hkwTHemngZE+e2hTwIeJ33d
3shh0AoEIPu2gU2YPP16MV8NAe7J2+ZbCOVfigsLOVawMKXXFdw66DLLHTADXLPXHffScDoRoncV
bA0MtfTX2KAO4dAry+s89LHaUrVryEp/RhrIfAb1JYjnLgDelyI8ZdeJBpWPoHMB0p1lHunlV+Ql
62/QAL6lU96cSbXj4pAmN58YlFnaO5LVw9tD7KsKkZT7gYNu8hNRkbTUl4hhwHd1r90ArXw1XeZD
P7nUUmrKpOs4EGRuhyYDlsZgg5+kMI4wDMbgStBchOxKIpr9ar4SC/c3+fIk4Qf/B8dABCR+2Gfh
clgnLmU8fd5sJbR//iRFMeVAKgmbwoAoWwg0awjfAIZXGoFtcDxZlgsQvQwWzXjahL+Lx+QnAvCt
Z2CU3OGIlO5LN8lbDMHuQKq2TOF3cP9N/ms9UE0f6DEuYmdTXR/QFxnFSrtg/cXmS0LQhwNrQJFc
+Mgf9oFDMQCK6UUbvn/g4dWtY/lcBQtemiM6Rsied0o66p3aFWZ8lT/+3/Og4ib/PO85wOuNu9uF
DpXL3TKl7uixl9uKnAkLVijweQaErgzVPYuF2mKi7Wupk8SEn2Reaz7XhO+OtelWZHAqoA7NLTIM
c3U6dpXKjS+7e1wJKGvoyrSqm+CQu5iwbN9jRqAVvpkvH2rPK++1kWdTsKgbEtMLe9jQ1INvmEn2
XFXlDWC427UOoM4ajG2YRn/oMTXCcV3zarfg7Zhe88TGtKZKJCOc14EJI6FONSqMfPMB9aEnE/1R
L8u+PUivGroFfcMUlnxsyIPJk7WAQjojxBjttGl15CfF/Ic+e3zjh4ljK72k1sW7DZ6kRbANOVF5
v4jU/t60pQxKhPdPb8aX/ORrt3OPvJDl4xwsWZ67JH5CRmQf1p8aKyamdUGwe6J5Mqp9soprgJtb
B1KK1xwn9DHetPAfpvICj1DsA99/Xb6jhn0cBhWhb3boO3f6nZw/i2OUU8HDguBcAcDf/lnZYhhx
MO9ySrxuQvnQBRcuKwjrH9phqKMOFgO/fcjfQgRLS+uZMzoheuMwXNxSFTAoS+TjY9zWjH78DNuL
jjUl9rSVWZ708NEVsZPmz5I3azNyzmTP5tBYHdeynpxp9emLtyvs2mMrOTyGuJzlX5NvV0bnwFM4
kkZ/WWAI9a54NnEmbaDqXJZrHi2v9TE7OMso7SaWVHjIksQPg2d4fMDcjMfH73+rJ/gIlvVBBiA2
3OTIOIc6u6MGpaNtP9cIijGlepuzH0NM+LSrkflDmvTpiNOO/2Zqlmw547cNtn5zx8u3D/n4gcfL
KUIPf7CU2BOTDOwustouKCyO34T4693E//8YX38XZcegv+uUduSTJReAPeNcikQz6ZvtPyISS9XL
bthLKJv6ALOU8yZ2lzqa0IMfvEUnsC1rD1mgsLfnqEyy23VvBZUAXeYalGYbqsxGmDjgDH1nA/z3
R86h0M3+diF4+Mu8NKoZ4HkTPjReAGY/UqRWJF3wLJBFEMwnwwpXqF6dj2Xrij7n3M5UnQt10Rgi
H60eLEYda9V+t6USZEr6fciMGdvmbCYvf7d3zDavdi8TRap1MlLnyADxfFCFblYRoCrF+XhodI0l
MoD/3uvSeZvQIAZtYruKb+dCDtKkdDPxAQnh3w5FoQ4GkXJzn3a/E+tM6FRwYLbDjwPErsbCzHWA
OZ9XClV2fmL3rm+6P2206eZ/cftMSOimJUsIw3Ew+x3Z9I9it0ZbvoPymDlEjKrS3h8h90x/6G9N
15jGadpeLvcA90twsENVwdq1JSXVfBc540Kjy0uVZSNNRJFSWmoCgGI/9c4LBWukJmaGEqEpKdBr
4FyJqt6bFHXiY5jogrZWrZbyK90H8j7x+PHhrey6RS1/MwW+3aoa+l+E1aRjHKJ3bod97bIIyXeW
Pp0VxMxOsSJfHDsFl7n8jdhYQVyTnEwJk2Johk6cSfDB/zW9FzRbvxptXhFbSTCFDbjRVp3h1ytz
FtejsjELFAwxcsJPwED7ZVh2zp1AWuWY7cw/jLphM9mUlbsReE6uuql/Gc4DqILmPm+U3EkcLKor
rws2DKYj4ge9Z8b09G3U27lTUyaGmHsGolNTTpEEcXBG13pd1WkM5FMicAyWv+E0r9It3Od1vcbb
GnVx3XnlcQsluDfF9o20/xFKUQ1FCx7yFQGb4jm8FjiKUIyXtTIcwrCEOtRnIayKrl8Cjd7YlBQm
dxawMR3EYsRxv+2MX33R6TTcmKR5bY+WkT8kg3/1xlBH+qg0Sm6Sswrku1xa6P8kuZpV3Zjzu+pS
UXEcYRwrQWXa16nCNclqM79tVFWUi3Fy7lCFHcC1OZbO2UgK0YypIKOM3tmU6yXlge/ds9ez2p8H
iKClpwlLbEiFBISa3IuAwWyj+1LXHX0RVe6VzLF3oPDDHoa8TEUYzk40foIcMMK6NAGSjE8nyN0p
/EK/sRLTbskv9fENJs6118gLeQ/EKjmreU4xvlyH4qAgAd9XYD56ZrRWN0tPTS3LvJTmLNJ+zV4V
PTJMjXTxJiK/xX8GXjctsSKG0EyYgpe7vR6UQXWM14V/p9pA/dPZqKRScFJm68rMnyfnataPzQPK
h0vN8uzZ8V/3wsL3eoccvLCmwQL2R+q8TAzryxo7r5nds083vZ+NVhkjf8TOqPAbqOk/bmXWEVWp
YcMZQT6Mlm1ceUjnXby07Eya8deNf/aIx6WD+ZfX9tQhmqPiFh2M1olK63kNo3nDsnoY67tb6Nyi
l0M16hMxfD4AkVSA9o5TskVE8ZB9ACqePh9Lwcz7S6kl6+ghJduYHbAeruTDK+JR2pPtApjbCkXm
+YE9k0rYX2KsN7zL3+lSUxhPYzdRxykyRmNoKqkyBmUU46WwrMUF8rNQ8xXn+9x+CCK4ShOxZEhX
BC9nH6Pl2RQgnVOFxZc8MAQImvvg1ad/INCCEVK5HkC+uL9F1vt0P0/BXYkqAItChcIMjI0svxtA
UZlfG7hl/4J342BiGj884F/KKyU4i+BxFtBPDwTxav3ZnBMKmfPcDC3bF9lXJJT60rzlaRglqh6/
Mxv4R9WJYERyRpB1WXdUP403WtaypOjMm2XEV3j/r9drGnolu9iBX8DTcIfiscyefz60nu0FVBn4
mlmg5e5CkdpBQgkB3ENqca5jJ/hn1AS4HjcB0hn+74mOpexH6Le+Rs9mVNt7l9L9Gj21P/8tZDGB
akqe59pUL7R8B5jpnPGTNMB6kmLR3aLyiT+t0ZSNwCs1R6y6wC4b3/ntiWZNF51Tvv3XbMkgRwnV
sc1EspHJd2+cIno9OYz/olQMthUvLw3R8G3U85+UT7KZRwwuQ/q0xzbboQg2J0wC9gAX5GxrdAfE
82OwHnACx3GyXBpsKowobicVvaRBJ3B/cLTjayoEjY6ZZUeca+h6Jy5ZwHmNF1t2yW3ha2hYEWIQ
zXPGtB4O1ZF3UqdVTG0kVSq9kudiz3NRmJksD5DBVb6JhNzNrIL6ytkbsB9k1HhrgX/SO1dXTVcp
F2p9guVyiShqZ1xBrTCsDX9XBAXouL9zgyffUhFLHKTnXH7QNNEcJxZK4lBN3LBrRhl+nl5ba1Eo
+UsOxgSEjvXs/i+694h4IjYB9PNOU52oW66xfrsABi4ShlfGx/xWjmY8vRTR17PeLgpZAtAlOWLI
eKA8uTIlA6eFZCWnleMxg3pZXZyRs5fakLUq28LTAJ4TXq7QSD8PiDU41uHvFvhxyPtkgEHhB9Qb
6Tu2paidrIEtfUc1koQxLHiKzynPNld4eg0HzC21nLKx1XongYMSQiLZU1Tgu6h7CJHul+LrQFmf
/vadEFDyvgxbombPv08L3LUxrWAabZtaiPRLRCUDOfp3/C4edQpAsndC/hNs41B+o4bkNmU4usSv
F3z2E2JImFL3NprHGn6UPOeCyzX72dcprmMubJV57OeZMLmVgDmfNeSErS64lP638abSS8mNU9sU
K0vhmhkDnIknc/X0d39eqAetohXG9TS2j4HnNn1d+Zw/w7C+zrVwZyLHz06GJOMTTsT0CWufnj9D
5wm4AHYw92HLUmq51i512R5bQU6EzbgLu1AUklTeR7d0Q/SaiSQ7Mul+5C9zz0hZau1ZjFFeV6Yt
NvZ+td6zbI4ZGp36T5tcxebaXxUGadC2sjNN11dr7lU19BosqayE4un9D5MvdNCXxT22ppiGljym
hDw79VMpaOVOjSyYOQHmEcakmuqZ+VdeX3uSERITLBiW+mphGY2BTGqoEYm1TJKy3kO/0g+URBvF
DnQdOp0eATaWY/xa3g2IYpcXgFmIS/Jp8t01BHjCc54MvqFqvoBWawK1yNsMIYvLbou1wVjazd4r
qjsRA4+XzVEVvYRINy+MPUntp+HVKecwsAm/37/pmMoHBJnOz6L4SGm4gK+9vCp5rAcvr4pIaplQ
yW9/luXs74NMzla0EjqtyyFMQrve0pfpM2FJKn8Q5yScUZ6gh3v1cj56KzNfeKkd/LNEHl6qdnTl
Zlhz8zjH2muYeAHz5hywDJGU0+dYQ+4G3BO2++BuScKtFAZe8Di3fh//J3JTj3IhOatCu6mY7Y8I
w1lbRYG3ySdTlNK4vOiv07C5E33bg/ke5rQcICEwa0o0CZIU2yqBBvW05u3kaRjazZrfvZR1Lr8a
p7gjBIOsWv/TuTQGSI71jvfPBRAzVokTux4m7sNU1Q+AZJMMd9F4ugCDR2OSFzld4XAu+dHgmTGx
+d5wYu6i5XJ3pWQC/pP1z+WEZ6S6JIRs911aEqj23QpEQsKKnsz+reK8/ihox98k8mGm1zHwq8wZ
g17s0KDxvQSGQmMD8WITqWKwbZs/CyhXy8amZxGWSQrRtlHVloBYoy6l3F8t3SW7yGOuI1ZT/L9t
xpdtMAOGBZegdi1zXlYs3B5cRR5LFzk7oo01haQ4kGZlxBbNPN322PfpQHwv/jEIsdeIBJBuJNDV
vTE2BUUmWvVBgxSb0LvQu5QPiz+M9HbaNVck2iu1riCSC0OgQ9oHPRl4uhZRtI8c6zKaAOMkDX9e
9nAcZx89eN6I6MRwOtIP6uptxqwsm+u4J+X2t+Am3ETAHm8Vu+GmePkRZcWBrUl36MlVimpyKQ5U
lARNfsn/tTc6R5QKoqg7PCkyrC7pzVL5FosO1H171SRaIQmYYla82FAyBimH9zJJ1NWc1KFRQ8J/
ZmDI6YvkXhaVpegm9Wpyk/s+/uKx4PZHcC6KNAvuCp+h7kOD9/nVmuYvMHf1a5lceSVH/ItWwFrO
6RPdM9WKS58RmmyC9Kh+nbugbxN/JpvljvVvCSu0F8Y/OoDxeq31tMtL7SfNZAUpRHzQBDXA3e4A
C56HIza09FG9DADOttVb9Tiv+HjpgoMQlLmQMRAUbV3OfVfSrOcUNWybGhCy1OMlX2ejaEwQs2ld
KkG9XRVb2VNdRBokj01QwA3CpRd97aaIMkg9he85PLf0Dqiz73Bq2nM2/cH/AKUva9JfNEVBsT7T
q4HR9TpTOFhhFTdXHyip8vV7m+x0U5pPiCdtPzoU2uOzVQFotngj5lSAYdNZKQPpOgUojpm5aj7U
6dHJXVfKBdRoplrbBrS/8svxPAZjZ8ZJk47Foeih+GnfuB5zz5BEt2A7MWw3rPHANiavyl1GM/kV
YrL3lKq9SZ+8dRMrFqmsB1WsAghBOxYxP5PGzd18tnWJ4QYobRrmYaesxApzGkdBuR0fncVGieQK
x83x2S2bp9DErfpm5j0pOuqdv+M33whnxK3VAUxdm5h/N6Tq0D81vixQIiT4VcbpCAv1c3kZQA+V
dYTxi7n6wDzMihE9EQm0XiiIYBHiJnf5bv5CwU7WNKse25j7aPIQOi4A7lWjN6otAEtNSirROub3
yxNE5fHFYbASm5KUeYlEC3cJcL298f4uH6V49Y2qzQl9ANE31w+F56+wzGyP2ufL+xybUR1DfBHH
xJBa28bo/jHdK7jY2QnL4KDa2L7W3zjb2tRvA5fccQCng4UBXPCUs2TrCdtISxfbE8ZGxCAP4ei9
Gl517YcnarHJhhiGfbBX4lHHkjwgAoc25Q6G4AVae2sapBDUNfZFL3Aewx9ptFyY/n/v6TSAXX0j
XbNV9/TypHB3xIpd9P6JaHSmpLBHc2LD1WfB77IubgHVw5faPDKq0TplCWHLgiSwM2YoZzb+KQV6
GWBEHzzDqBHqy2KLwt0I6CyFPM7VI9oyhBAbZ4nVRisXzsPmODaYmGJPok3BuevbxGw+DPLorpvX
uP2gPekH1oEn7KMRJjbv8n0nGjIaLamtQHWuwxtL/EXNQxp7gLru0E78cjUOi1kN5cxQVQYFG5d0
dlkVXGyGZf4T/MA1X0ytJuiujRgjusFZeiueOF1n93h5UQ24TMAE0eomySnFVnr49I+u3Lkfl6UL
3qs7fEnsTawJZzCLqgMgO1X87oSM91TE+IuapbSmsrSbBBBveUm7880zmL62Rg7MF19mBBnC+ZVH
DEdKlhWpBSmFUzAsXEV4//4MsipM5SUYlcb48vLuH8SthzZlS6l07lKvjNGILMusxYPE+WllCaB8
YKlhQGTfDJpXBsSjdCWsSOyWCk3EDYKDZQXnXpQiXOudujXxQgKjpJOcwkLa2XmZuITq5vtHWayl
p8i7Eyss4Imsq8qRIkVba3Xm/2/BUOpAKBmBP59Ri4yS1N62z7Rk6BMWcmFak5ispD90M7UPBmbJ
gQ80YGmANaJ6n8qTVN0VIdckc+gq4wq9QE52ifmT7uY/PycN60twXgZgBVbD7dRPtuBPf1m5YZNM
e+Khjj5kN+TSDPi2y+P1nvTcy8HTgP4EsSACpX52liWgEMjDnZDe5MCja8Qs2Tc4zoqtpAE1b0FZ
x+7A9Y5PBFlwfBSynV8PNYV4H5vtSjVlRbchTMx0gTFYMQvPSmtFiMRxpZ2bzSfAYPfSLN2nYtTD
BLJY/HGZar/juF4BOjIlgaRsbbvGnoH8lLivU0zmfgq+EpE4CR1ol5DtjXWWowrGKh9+cXGErgev
0F4gxsnwG3IuT6VV3GtALHUA2xuWU4I50zMPMdUQZgCkZicDnvrgAsoL55JdTIKXer+ygA7m+UJ9
ML6YMnPpag8DFsC0IEmzXXVSoh24qf/mnw2bLG8VSAwbZ8fiugzXREZ0zJkev2SqzFS/6Y0UsMJu
6uXrb8yNgHIWFUWnZ+mK+3GC10cVcBE+vWijt6LOFYF4kmTI1tdtsMmuZClmY+5OmQqd2peiBzFr
hbaZU+Qt5nCs2a0Ot434vvphc1NZRey6JPpauUHvObsJ4C7SY3lEyPGwhagJ6Bdq+xU3S9TiuLT/
+aORN/CgyW7kZrk4rIm/NN53zx44KiLpPrQBh9UnS2GLrUpU8zR5yStZt6ApolENpPZNeiFhWEn+
QsosFsPs9pAr9AcGaTjOjGbcBRXdII4ikrQtXqad5EZKsD7o+UF9/pSho3+9V/78p4jmJz1pV85U
vOX0fJ0Rns2XrpLEscOPYVn0rJ51lIg/LuQneGSHjulvERGlB3Q2dhdRLs8MA9jWKOS8daEB4csr
bjgKJV6ATauk4vhplS6YPPS4k/QqdvTrt93XGpi4S5Er2uU2rQ6Z5eudIXnX96kniLXoR/nXpSNQ
Gzy1w3cHDDnQ0N6Crvv2DvubclgR004ro7lpDbJkOI7yVHoO9fknY25wV4YKpYe2BhmB69Ma7BX9
njxh0Eyzc12A8b0b5wzn4/hGsAjRgHRgq0blVu6ZPx4ZM7fkQP7DSnOM7xGDLO00fCG0l+NUtuzU
R4/s3aCK6hflI0gX48jQJ55j9jCoKghiTPaQ4O1xKhR/LgnHIHfcz2du9HdvBrZvMEv17lQYQZVz
psi85iSA1Vo6fGQuwtKtD3coa9eQUNe/AR2OrhRSShGwzI4EEI5iVcNTYmZSs2lOQKBPl49r0q/5
ZSZs96joHPinUvT5g/9uTcD/XXWWzVHkgjyEYUexQOg4w0A4oyrNM1aexuf60ZKhjCb6KD3B2DsI
aoGHQb67oxQ/xme1TSY9dY2teKqKOg2GfF5DYZalVZ2Pm1Sw7fMNd+I3K2tNdhOufKi62BTdMICe
pb9WTSFkL05acwKpxW/DpMkGGKN4AZXuPS91dyCyDW8V8Gg62Ac/tWhEzr5wTTDSBOHo1QE5Klq3
HFgt2iGw6Ut0tYu3/bdcZczu2oaW0qp9yy1lyTZybcZbaL9FrG1zHvVlHhN5qFfi4i7IowFLibRY
AH6zLfeL79C1sdnWqpy5X02ICk3+sub3NkprzKoT6sXOgKKNadC08mEJBhWXXmtKc8Xb4ke55hpu
8dB4jEtNAORwU+4RJJhe7Mp40If6mlmX/PJdyZxbQ1EsL+ofPAoVHLhw8NWlVKypLl7IwcxwpL1g
CyIaQE4wc44htfjcywKBWOfxF3rDngY2upRQCEcE8IwOyTsMtrr4JDFGoHfh9iiXsHN0T5o8baGz
Mz0q7usCLntc3xFAbzUYSOjhi3WpUVrK+ofbxNtSX99DSGtDxDXP59LEl47oRvFmQm3Dk4LTv2YP
/8FAFOObOgc4217whvHLixGkwUiXbJrR4erPk0I4Mt/Qfyo1XtAeyJyh068GSjCIKdRDECFzXn7G
73Xuhz4Zzr7cuFbJS+oMJT1FQwA8zWTeXVdWxSpsiDzZWNiHidWuMJfyFuMueprtDE95HPFlF19G
aqRKvgtr2zkHrgIAvDZXcAl66xXxg+3SVAfC08fyjLlecvlscKA39OBtjOrhiTG2U/mg16ytZuPn
J4xLA9Zh7Z30+R1UMNWhvOsE3nCYSrN6ik8eioOwrBg1+IHOD2RLbek4JqSBdAuvXPNW1AV7ZUVr
++vty/FDU6ZlrALoKpflDectN6rdqzOxSVB65jEJmuVY3HDqhmteozn4Q6rGMxCUCv3PA+g42KT+
GVJMlLexmXdIEqqosDzHf7LibMkkfeKhKGa1FaIX8uf9QbGY23opCp45N7pKiK7dMjZfsLRYzrKj
HfLt+ljD8ieEOo06FgdIZMjAhDAcl3miKJRO9J19aZM8nTi+U5LMrsXObtq/kJlowET6u7cbv4m8
NAuwk70qZ8arW4PJDUa72rai4sYpmnJ6qG5NZofEXYM7cOGJsU/t6zXZiPA9GpJl+xNJvJPLt08m
782GjlkjGvuGoBbPBmYzNsT5pNbx2wlRan5UNHwFJ80bwjI5xnNjJZk/g+9BqlaG9v+DAxCTbDKe
raJ9wc1XOL8tUt9BWTLmmptg/GQzgLsDqcZGJrAyeGyZx4E0GGiUKBFRepT6tRowQr9JRf0JH6Eb
yDbr6fa9lV7vQ3lwOvxJ7Qc+G01Wp3CGVVKnsnyYcBBhZeGZaYyc9LQNguhlvkJo9dIn7FUucRZo
di3hfA7dUUZmr4+Uns7TT7+nupm3Vd0GBXBm7/S9FF6t5xogzJdqBdgXKqWbYvwPiRtrcsWS1heW
nKZBdt4E9gVawbUf6fuesbdUK72qE4DgKRX5mAuP4pGpcB9GMYMFW0ifjePpgXs+2N11Wdn8GeII
sepIr2S2WJjeGnI/3zLBAhhz5Or/krcHM38TgQL/e61fAg2mqQ4MC819AjNwOyWQ0bAdUjeSdYU3
zYOG8XRfeIaWK+wFi3JUVnU8kVO9ps0joBjSFiY+3OTKpTesT/ZgWNXgp9GQI/ZXGF8/3NFTZkEC
cDs77+febvzxl4DrZ2UWw+yOT7Dp4M6KY6S6+eBqrxpZKJHe9T2/tBLeAShCn/ccG7RRm+slE7Uk
TQM7s0sjZoIcM/UQtYRNanKwv0jVUmNQb2tPNA1nzqTL7NhWhHyHlxaD8TDUQb1FGfscA8UEApdi
ZfMXs5kGWY5tFo/Ihdule6QaUOOs5R0a8qtrWPbN3xQZS+3ouwAHjuQpnWCSHjju+zmarKCiMKgY
UdqOfC+RQtvjuFqeiiPpaMp0/M0wVWFBgGjRwt5H4zb4T0b5AJfe2Rp5pnkBySTsg+BOeAXz80XV
q5k7ekjeDeXTv8IJbrQxI741e0viSwA3Ebn9NakDMKw4cCt3fQHVcJ8YRVUcwRXQkFMZUbpZHQ1T
el7/KKotpHkSerzMbQdUtYF9j0i24e48bq4SrEWVPs8k+ExLGcKRWda3e6uLTZJLQs/4dHpNeDmf
Pc1R2kfqp8UceR8LabEcm5JR2mFcyUmpLclkg9w3oTBgrxOetXgUa6FUu5f5nIJWJI7CUqlawN31
OlwFvvsU1LeA8IDAFNkDoJ/awldDumcSTAuH7nhaLY8uKT4CKF8XKoIaTCVE4ByA8gh/vdGG5K31
827SnMp83AfP2iktOqITKDm3R9zoYA860s3hi0aGm05eP1gj79MbX4+a7YAwtZSR/zczjhxVvBQO
6XGgWbza6yTRDGpOMZflc5WJX9HciqUi0REkDEPeCLlRRHSFTk615hE1FC404jCPejIubYCzMN3z
W/oOMhoTfYOjQOU4T58NUUYI/An6RWAykWo28lX67JUBPqyNElprzBf9vzqDSIM/9n7WehP3y8T4
/OpaS/NVUJeGSQw+MdMl9IOW0t0aTmIYvgwKSLmbvj4+DST9eBKsQUBahQ1Rx6hAvCSgIB+NKf2k
YbsHHEu+BEpE8c7bI9sZW4Gob5AouWdNZjCT/k+cCPVcCvHDcBBdsUUh4+P4N+XJOTZNmTtGNIG9
H9rLh3i14gnoD+IOJ7IFnkhbrgvuOulmhdI20yB2zy6HDgdcIgtPVyhYkfkNUci2kMCOQyWkhJzF
MSi2mokSyWwzgkxSu0dG6EFS1saS9GO8oeL/Z/DIsKVOE5yOUN2QFyE6KpaoodG3xXKbCgPxIQi6
sE0CnRFMVkDtYWYGvbZc3PD+bgxTgL3oKfW6ROf6NTh97OwcLdbBFMjfVLgF0OE0UyYqmeeLry6G
4OPImNehNY7exF622B4QSB9GiC3c17ntbQbSaUFvP7mmtSHj4wbedIRwFu+gKSMcZ4Y8jnO77EQ+
BzkbA3YuxwYrpQUZv7jHykQaH42nFz2p9SIlMts9Bdqexgaf6Leua5EnE96vRjfMHDesKxbk/M5X
YDzSZenQliyUBtSpu560wTfpHsx/jRbd/n0+59fBl7Zgsl2tXOar394NtrLzElCQ0DbzajgOmbNc
Iiq1upQuu5HvQ0CXuRjCFuLa68eJHrhWHlz40byx/LD4kI3XxcAwRs9wCIfnwkw1wd0gY7/ikSrV
CiRsv62l/QGVFpBTX/xnoV6wmFEz4jDFkjBt/RydMDSluFWS6AwswpzAnfeNDqQBEb3wYP6aPHdP
RBW2jWExFLpFvSJA7tAh9KqzrRXDhFRn0Nn92g6/2XkL4hNa0I+SIh7jIsynToE/aYpNqoOkkvs2
CW4zn872Sq2rxxHTfX1h1vofYx12tEVRpS/ITU4+003fmx9EorJNr0IqHSyIpUu+9USGbuXtfNAh
/7tWF+ibtXTGuSH3/3eE9cDba4f60CPGz7PQ7bBa4HZTq+HRLgecUBnEebBwmdZ3UVDUaD4d4yLG
OG4LwBwLcMgYG2vgESW3U9gPd/7fQ0vpEecuQnmFs8HJkv82m3b2MCVj2xXchc4J+xfqK9UG2/4z
JfCTC2yjXMm1vtcU88WfMh6f45VvSv2EK8OmMysKujUCxUsui8Kixni1PXk8+ypBvyg1mhDxAGkU
myKfrOAQagAl/KmS5GaKoTdk3wDFbFkkaZxxWDkIky1fS3Z9rRXvv4jus+pW6x0IDniDL7YJy3n5
BqK9lWt7XQf6gtk3wKZonq/Cc3uRFRpOfESyJaiL1IwoKXH5e35xhOJ44zA3h4FhD7K4ileUQFZa
TIFiU+ZOle0VzllGTZbYx42tPTgiocoSLOTwymNR9YCs+mC2b9/QmkRSsNslvM+9liwACo2DMBy1
X5hefubKsoJJe5cLCVl28i6Fk/8u58JWGWQnqScIw8E6DYgRVYt5KtCTkTS3JkVdx7BbteUTRJ9d
c7gN/YzqR06EpDhJtQhtG37KW5IQMjB/09wX3vJAvOAx287BNiKWXRPRFssyoWOhho4o0hk5cj3R
XMRWe+8jtz4CLSDmJl0PCZqq1Jq+Ab+u1rmRcrrFqAXtTiEONvYVEEkqLJ0jgYz9+KhvJSWTNcMw
I/YWy0AbkShz+/vslzuwifuGNQ2ck60NO9mQ5T4CUX6ge8Vtxs2/rf4QJkseBwly0htl1MDvZOxS
HEZMrPb5xfA86d1LrsPFcjkJHRW/Xr40rR96Ra20h4TVmyDSVjgnRA+UR89/gf38dZuwqo55YG9a
z66SmSFgrqHsk6nn7iVjv7/btSK9jxqo4FVQ7K5z1681YVeRQAygKKKYhL+dsddVeyhFKWJ+xdjM
ZLY9PR3Pn4a6cGLVCCfUc/uQOxSHyGzz+tUWw6Ud6SMf9hEqkrZVzjFInREe4oL8JVcDmmW1/+ib
WqMCdMj6DUjYGEjMdFu4wE4ujFsE8WImzAP7z9Ho8iI9X7m5xtB2beMSQ2xieG5Ieitwpulk1L/K
7xPOeMWonK97HsBUhM+lW3HaFnw9RpypBLPqzN/u1e4EqRclnpyPKyGrl8VuaRnGaBphsGDpO/2R
YDgKRkEBMdK1DDaXsR9nR5eQHlISt1uknNGjfZKciQE7O+Tvbsxbx4PtzXoEQA0vRgLWPIr1j2gd
vTkYCiL6Ky4/jj/H8BPKi65kVudgd2sqawKkNQsu5rkBJQjtY8uTVA53Ccr1S3OD3eOGY5tTEK8I
jEF9/ZD0cBtMflYs9PW1c1KnzEWd5gNICpav6+cWoqEBmXUE3DpzZ6VxIL4ge5G77rC7gn7TA6Xv
xa26ovVTGAifGU+vvfucj99B1q01hCAVQ99qfsJeg8QjIJM/TZV49xl2q+XTp4KuuFZksacpawnP
sZfrEQ1WisSwekctKGs3pOtooE07SWiWqVmzE7HCYOJRQmS7RVB8I+tc6nSROX9V9vdBVA6N6CZt
Ggidig0laUCxzL2DLQRmdHfXL0d3fLiosl7+b/Ym4H5qWtYNldWv3Cpap3lOvSDTZpaGI51oxX/i
edgIdjrck82uoYxfILpKZHS7pa9pafaRJBJh5xvQrGCwXm7XV/R5mrxxnwG6oCPzzY1SVcbqD8cD
JIfo11ZqfLlhIBRH4NErp03IURR5Ih9mhPBJO6daJ9NKaGhaSTSftJMHpAxzMctBck4+E9Yz5XmJ
ZWd2nZrEsMmA5GZZ1UuF73AhAQGUAJRqW9Ds/L9GSz4RBhAHkioMLMH/7yDc49X/0IxikqEAISqd
rSaZXoNfGoFRLjkT2yvKiln062BmLZLjYNxGgz1oejIpDG5lpO0NDB0/rUZKFO6mQ6RqfaM2TTYl
axTmV4CkoQzgBE9XfmGe/xlNxUIpKvk5pTl0Bs/dMHv2/FcFJh36+X8paF8+DVoG+WuTJEZAWosp
7elj+c470F9gjPENxGLCW8q9/R1jVHTORim1dUZfVAy4uFHQRPBxT9YQhBDKkxjk92xY0CeFimb1
ZEyf/39qNMUyTIG2f9ASvJvSPZQpbDBMtKmM1M5BwW9B3ljAoEaMq3egOl7fZElyqW226GZi53+8
r7npbUjKqwdkVxv2EXbTqZBDjHTwMpHUcj/C54Empd+UN8H06LoZiQQbbvietf7KjqER+MG4zKcQ
T32ka16PYQFVj1ShL86yG7nOFo3FMLwao2uj9nRCuSGlzXZs2iQbUfSGhuPlR+4rBcWfrHMCiq7V
HIEfU5S6evulFYLDLF9JuCC2NJxEJMkQqMqA/dRj/YI77h7Jbyn+3z8ysuD/Z/xN/gSYwX/JZIzY
kS72xwRp5mU6GxhHoX3q4qOIio33jaXwE2Gt/KZwNo0Q6NTtwNJPuxgk5S84opi7g22f0IGViH3B
vJAaspTvjixOCnpuWCGs+ukODS0kAOLY23d0+CMigQqe+rTXeXqhjg9zVlmSx+oPKJ8Lvjvm7rnD
VbhzFOVgP1V1eDtoxptoO9o+6X1bYO3K7v8GT8xOj0HmlTcUg9GAJtPun1cE5Qwu6bwxxWLDfjRV
srP/TVattWe1EkOPsoz4nYsBZI3ELWb8rpRlHDP4MYSRPdyzX/rt67HjiLGY2vLBwOQwAJRvw67u
tQjU8g5MSDUP17zuhCeAYATcOaZw0/sjnhhYlMgWRT0/2ZKi36TTEPpuPyUcnxRALB2uCRv6zcnz
iwhAm76zz0W6o0ay7q2ZG8r0KyV/GtWxB9YX27hKtgCYMOY9x8ymX4iJxZcBh7DPm97ahXcNd4Rz
AbamK5FqQ+V2H4kUKPsETrvDuDe/dc8huRTmaFi5BU0le1G+h14JCrTrC0xkPh52v0kidmzRCIjx
bbcpDbp3H5wOmQkF2uJz4z602jByT2haHFNwqp7spAiVuDQXS/NI42F2FC6yPdfLlslAiXiRxCWg
PTwp9uCE916UU3S8/VhB0uhPsB7r/2wv/cbOObZ/etoVvP3WIRw3yTJY1cjKkH26Iy6ozx1pOhWt
x092gD35nleRtDSXVBmMkr5f32vteSBu5r4p/X5tYEsLDvmrd69JnlEyYI7G5X96nWeYJeVudpCa
bL1yDzRmpW/EZCCA66NfZTYBKOHs/FBZgm+6h3rjlihI7odrp6CDRd7qH6u9KJOvV9eLNxRfz1yG
aGM/a/ehbSE8ar6Y8e/ighQZYvVXReIXHd2bUFS1gfitHYn3ktp7ZqOJtVrbcA2bA4p+rUlgvJta
fi9KWClKAzo8hBHuFTBxD0WZAiryiqxbhRlu5yztLe2RKb49eJK2Nx7vNo8Hl+I/aIVdywSQa8nE
9d6WorOvhnb8i0tPteez3klFtxOaYt0i+eOQR2X5wymxnxGbC4BZTxjRFyo/Pbcu+u5yjtwe8Xyx
qY1FM1+LrD56Rxg5J63J9Ckr0mCcY3/0+GV3t/s/j+1fYzDKt8cVRDC+b4yt3N/ZiUBsBz0Tyvs5
Ob5zGVyj4xaUu2KwZ1gMvQlj1JDHfyqs01clcRTEINa6b4GL4Me6cYjrNctkmju3WDo+h2vGB9Oz
hQzz8uBYmuWGK6OOwl6SihgJHP2vXcXBpNzjTMAHEVsvk17GtXi0tdcapnoxI6l3a3r/kGV5E+6s
I4X2GDUm3EvjoPnCIowtGyZ77ipXwpxe7pIyaR+N+lmROoQ7K9HHe0CWv6un7+mvEsIJR0UQYY1q
ZxTAjb2UfROh62hXwImBcep9DnXF5WKt8gC10ILtr+MYil40t+WdPuserYdyNYDmmmH37l5dS2CK
iVJzzE406mMa0CSPJoUN4jyZ8ehPWGSgsZOXOEhron2Kn35+P9e8aYviArONq9jYsr3IaibXXqKp
Ggitf+ldHZBowoEp0fRo6gJP6WUKyyq34Ob/H6W7RwiWHHXo+DKHBR3rBKBKfxz7EiZJMBcvA7XV
1HqG4RhyHjGLYdEf/DOtCYzBeM5kwsIpUwy5kdgCDfta+8TceMH8yaWjaPaPKUQo0Sy3KwyNTE8M
4F0GI0HDcO1GC1OacSTnQqdb6e7hM5TxCIME7t2j6NrFgI4lrOZ0P3NereWtmdIfF74Dh1X5W8Up
nTiYw6sMoG+sA/bTyqX44TiC9/ych3xJbYjZ29FoCEreNIxI0tiK4nPsYfXfI3y5g/pSUjbkq9xX
iiji1rm6mYENUXePFsZtilX9/rPmxiJ2Av0rHZ0qGc+tVSz1g4+2HfojCnr2nIX23ieYk9Lp07sJ
Y+KL1sIdcknfRcuXggSNRNWOxN9NBBJKzajBjsuL5tyhmTa0fGMtJZvIETefPoTF0UfUZs1ef1/q
AMtRsy9Mv2ahOiluYnjd9ALmws9RpJ8A9tQ53rbdgjmTk7foL1dqv3ZnkpRh9LMuH0cWDOupCuyX
d2Nrn6Rwjzr4PPzxm+XpVLKnXyr/TK8P87IllmjC11h/yo5VyoAqEi8sesI6t507LU1XRLtzBr3A
MRx/xRoZdIkwUhP2zxVjylp7oyOA4E/ncKj5PTigjAFr01d2fpI14JiAwtSkPBHOqyPDSoADyF/C
Wh002aqk6CZmmoAIDuUMsbhECEwcK2IA6siSDQgaqSek3wMb1wef7zqkRIY5Smm/CnIDTU29wF08
zY2wOMsH8lIlwRNO3I2m0byNKNIBuPrKpFAya53oELnHUsTzM8j8wetIdYis7Ppd13KJAuYve6Vg
nc27JiHG+CwBzt+FgfS37oVfnBgFCkGvZ8LnZ1zm8TNP2G1y2dh/LaqqGGans+BpxzK5yrXJZMku
zCjHWO9f/IRY/betBP7jBBKuaDlVoSsvmNtEjb6h0g/9k39lUoj6U7hMg5fKJCCh+yYEcjxmEgX4
zwto3DnT8/97Ab+SJF8XmHP3o6y8U1hF5GzI0Lzp5suyD1j/WIo8PecZOAJg/IPqr5AFbMJbZG8I
lzo+glvumMkHDByY66jdD/1DjoQQgcFwfNmzluxLDOwKBzNpP6f5c6JoRoQj3Qa88eQnDMnijc+k
vj2G3CRgXLten60VvoLjhyc4x2jNjenslFxJ0ZdfTU+c8H5cLQkX7yWw1TtYI1X7rX2AfVlWX9WL
kep07KmV1v4CvZakx36AnkziYwLnvznT7un0uIwokVvoC6ksk7kPLXV7ZFvI33LHXYWLXonKeJA2
vSgOvFBzQ80t5FZir1ABRyhCsjzxlM5RFHwztwsu4B//HMEpO0+tIyLummQYnY88RllBxjcjV9vg
tyeXUFUMEF84RZzHMQqC6NPNvOL8/EjkYH7mFCdvTilTXoeBJqTMm2Nm3bp0zpXD2BKFC65OwGbY
PFsO16o0oUqZcbsDBSVWkS55fznsgmeocaX1BrV7NDCKjMih/LTN4iOXd5ZVqBACaoPV9PCQVj8b
bJm1j/aAIWIw/J6fl6s1bKPlweGOMgqbmiIuHij8COYANJz0oli3xQDCImqPSXB16Z4b4mSrMWFN
h3dGtQiJU5B9u5Em5TL1Q2Jk5y5cD4WzJkwLgF4UEC0OLyWmSIDhvUbMq+ymk7UefDkVNGNzOKW5
f6Dq7dazYJYrMmFeYZqlzW9Ok2E30abi2vleV4UCSpR94tqoy2BQvf0Q/eOqK2m4XcZqURwqgAsa
Qt9+ZM2Gn+QzoRMZfzV/Vt9sgoSqx02flinKYwF2UC0JIryAOnKMzKLHk0RrJN8vlRcFEFSK8qFx
v88lD9AOuxeCFRcgR9/37Ado5P306O6CUtblfliJqq437JuUjGA+e6R+MNEKDJkkTNpZmTiMx/nn
UbVXuV2+PhL5W0stIqjwIdC8rDxadl4NNN1YZRsuLPJnvgJfaU0aoy2Ajt3Q2KD/uKZwVGI6Weps
oftDKS+beVMrCDvc1yhvjF21chBI1cmqdvG61UFWVK0i2qsfk7/3tEIATat7FZpDcbivm5iZh23f
aHKw/NEiIwBuYlRN5q3+96wMcu4QKQc5EOqsGnylL6LxeP1ZBeuqlFNTZms2g1TC2nbtCCcwNCyW
IbNk/TEFrbaISKRTxa7uiQ8nHE7Bj5dhv9UM7yEYAIGpUu/r+sV7zpoEuWpTMkwP1gv6HDK2s5/6
WVQzcM8HwLmcu53lftponX9B4Tk33RWcvcjd3w1Q0nr0PEy6jMFivmsy2iDkrL/I4xYZ1DOtgmS5
jD/MUqdT4ee9Vk8HNRZT/B0ZIVT0L1q58y6X5V2h1WBYlWNaUvYs3Ov+EfDaelwyyv4tkJQ8D5I4
GYlBLIOL5WyAFLjxMnWEF7E2xRfKu8kwutw9etr7aAi6d3qMiUZbF8KjBeNpWgJ4G+cSYz/tbns2
XIKnwO1AxOPqRWISiUN4Gc73AsQ1RCgFGVTJ5seRKB3mlLmkQ8rFQHJcc9fj5eqKmQIygITMZcuO
nMtICven+Qta5S0eM/0/NUnudQV/cIY5pePGTN0RGIAimnJDKjFzxUcBj56jQiCiMF1rLB6TuuQ+
tAszMqPqOae0CO4cb92l9wI00+3WMrBiTma7ipDG81aqoLZX7eHJ1n8jro4Qasu8j/v3rNNXYH2B
gK/GDm1b5PLvNLxzPz8JNSG6Nxr9kNffT+DpqvzzzR0ayr5A2UHnGt5pzaelaAwzcXFbYq63ku2N
qic+gria01TuuKM66cRRfIbdRzYWa80T28OHl/7+CvOAjx+fhymHU39NsAUWcbA7OHZQr8ymGap4
fOL/3Mx3k+dTouVdzURfwdVIGvXTDdsGdc5zBwo7duLdKC+I4WZGhqHi7MvPIisR1EfV9Y0Q0U9G
sgWqnsUAwIFqmwCZVcmvG3uOUilbVuRbd8dh/8MVjEdgGcQUa1K7ALqmQXiCbhrNAhq11IsqxDPo
jVM1LKiQS+PeBF34gCIQewAi2Vk1byJbHUBwlfjrMyhjuL6v9+7nCIMArrme1JCbmvtDitKic/i6
FySzCZFPeSh2ZaZrSx61wb5vhwmUCccSC3pqn1G3IKwTGC5xiSyBlpGzRQfo1Yt3mywcWv1+wVfl
ukkueIJR4AEMzRpKRSx8rRaf4hjax9gWePh/5o7pU+C5qoTB8eb6X5lXarmFHHE+GILFRQ7drg9q
Ww0OeFPkNGgPayFzN5eelZaV8oApviZgiGpMvlsegixox4CxSDMLc+Mq5IlqyFTOoDsYQKo1J8rS
buiLo1kATf+61HzsJY+wQCYXrnmRhf+6zSl1CuoepFSw7CEqah2pLFJT3FkJCSN/Mi9Pk5M/8KNL
5JAuZqI/nr7AO7HXOuEyttnSIUBFVUScJoh63X3SGNxKRY2siIj37OpgGTTmNRzaP3vRzoS+3x24
x/6W8AbJ6NUKEmCk97W0WnnFaf/woWzckrZXo/KAOdTWV8PSIQkmy+wvn+dP2CjMD2tcclMpsnrb
fbJ1hYiuJD0QsE5oQNeqdd0Ob5H3NDJwrOWm5PrU1UfDdRvPHbDYweyjEIqVzpKDeO31hBVLWApb
vYnzegOPT5IE2g2xgwS2alahHvU8JBgXhjfNlV8RW8DWvyOW5/DCdyqlMOl0hbK57PaEthpo9nHE
3MbmwNOPEEYeauV5ZFu1oE3DPD1PW36utVAD2r2rIzMBtowTefKeNkgRpmza09hforNZmwLXbGSF
JxeUdaAkxCTZG/RQQchKSuWThxZHHC+z8ZLnGJXPvKif/fDoskCA8HdOmp4KiW/aRUdhkbJmsyFx
P9W1YNAsyP7KvCTeHPcPJhITloX3bILyrESUuzJugkhLeSSqDiyd8dAnQn2JEKrtGoHSnGxNeZjy
R+Wc5co1vYmr7zkbR2Fy6bM/RDcL/c5EHUPEGlJU0X2ITZrKT4ZTG2Uaysvx5fcO4CWLbDyoubv/
MsBdrojuBD5DMI8o1lHdlOXem9j3csAXxY03Pnf0+DCQ8Vrzhwet+/aAws2BZZ8HWhjHbMKkcjnL
/dfW0LH78OMs9J+yCjxanY7nVpAAwQSrVKPj3WK0b7HjYLg2cnAmlLnYjlR0EvztFRDtTwJxq346
ZAHEneoh5Tb+3mGc6h/tW9WsjgnPiJNHhgvLcQ1zi2d1skpQ95v63TDTcviAX6NFmEqB6Z6JG3if
uqQn/z7RXK/2AlDeOz0nz5HMVo/ivqpTGSJr2TiFWtmv4KcpRlGj4k98nDp7uu3lo6He44bhD5Cu
9hn5AcvPRoj/EfcoJVfkg+D5Lt7L5zZkibnCalNxoiIQEzbGoweMv+EG+/HUG4Wy1DWtaPRZp1mA
xpzaWSNvABDD2j2mg/KbLEU1G3eEa+l3+czTOAuwx7R7TmtTX4X3NAjgWjyP+4g81pA9qAVZY4y1
YjUS6Fo5aEz7yWGF1RnEeMTwERQLOk0Sem7kmTOMpTryo8r6BITa9/AK+aPasIJq9wkCS4MCa58z
T7wLpItS4Uet66S/VNZZFU+b2pjtywVrZAfMeNKrRczKxgEYJwyiBMeyFGHCVIC9225DdBxy+cn1
lV/kEp6UFBcTs9izJY882vQEy5P/HsyZ88BbPcI4ypxDkOYEPBoggjjnBInir55nqOucRPTagyWB
EHSUjJ+ooIWl4r4NN713LranuVflck3Obd+ZOimVe0hUoOAmhOH9faagfhhCVghRZp6JGNDD/Fy1
Zp0Smqxrkwf4hfixCNpKaSqp/b5X8XvR4v4XyEJEK49IQPJkw5Mfut9Hwd0E5DArl0+yUYJQhHr2
Csa/7fpMtAOE+PH1r8rYp7A74lgkkI8xeDwbexAUYeBlPzEpGmIHMMXJSTMLWuZmv6AMOo08mF1/
2fZTLPjrXvMHCbU3hFvaWy7HHCerF6a7dghmCvu9epGuXgCooeOflS6y7FSzcOYlrrrnkQdJna7S
b1TytWVwHLYhS8/v/nXb4kh7pCqTYUu/vgB6WLfUvMUO4YK75CvZ0Z0i7ZMz4yPGEHH1omcSXeLC
sce6eL0iWGQLrq+imC96Da8d2eB9kzYima+k/VUwMnfj8WXlPGmzydiP+MdtJeWqVdTukV7Jea5o
vFNp0gGlEdLiHC5NSdXMbrOmKJgmSWKLflmORvu7RtoREvt5qBHQfLwwgi9idyI9uk+YzxvMah47
K7arF24XoLprWYL5YNLoGCsarDrySinpiBdIN2w+yYzlZpcCQ3IbVfTBi1IbcmsntQpmGkthpoU0
3qJjxsfyFnSLgTBkdztMPVCCR1t2PYlQkLVO+cOeKVCLnfSFyXyS3UMsr9m1tlPNHlqI4k1gPgUJ
rpF9Q+QzMB9cMa09dpkK+17nykYy1O6mo+SMzDDxMFNCrm78u0dYW90xmvk0wnJRgR9E9m3jLZea
v5ZiQ6um0w7bKIjHLUThi/dyH0vLG5uzs3QHa3qPbK+HS0ddn4VYSHA66XcCeUxK/rCSuEFLFZ3w
Wjy69uhWbpUfSzlMoKq/dwXeoTEedGAGagSBUCzwMKXTuO/j3DDjwUIQ9OHl0LO2QwRwmMLyIQTc
WGXNr2Gu+dSBLaLlNg0K6WUPGa3cQcqJk2rlYAWeW66O2dwIv0OEfwpoT/qIpdfOw6hOrFpzgorV
ALYAWPof8Zg69hm/7sa4Up+MEpJLVDfjJScPFGOEPjDVm9b+L4VI+12WqnKd4u85o49BGi4o/6dw
a+ZjZn/xpNrj0QZPJN2d6Eq0nMNDP6pirRUcgIIoMuxfakFxOZGeIQXkSRbG5nBQ5cuM60bWkTlA
olTwerxvyU/+0Mv/8mqDcoRkvM9dSG7SlrzmC0KTtumn70zenJZLMTBYSkOmI6oP1J6b/Dzki9uD
a1h2shoAepqK37eGOHdEX1/BQucz0EUAtCUuXIeUyyaWUVebG7XXVaur2zcnsocqf/F70pW3H2/R
VIbt5WjodZWLbShh0rAdW7o0QOyk5xOAooqjRMWVNZBIVHcQPtKhxUjTJ8sGaiMSE4UQm0cwR2q7
GB58LDtb7OV4UZKn10w9bR3tJp8fRR1AR4iRtB0/jpW5UdpuGu/iOTx5clxnRR1+TEgWQGzFjK31
NSafn0EMdPFJqoBTXAeb1XT/s3ZqJDEEqP5fWRLMoHT51GpMh8DvNYzUOFftueFjLzdYjEyctQ50
fReOn9726feisDDRzhPYpC8VOzqbdhD/JeuCvIjwkaTgd4NClUxTz3Q3cPgZ5Vj6C9bAC3k65bz9
GnCFCOP8zCvZYJJzyWuWjCL8IcCt1F8GXuh++y2ymmC/VZZxXIWbFDTgB8kZ5QpI/u+OR0Gu8tZH
jEZlwoR2GVo6c6zUa7SpL4zjDXCl/QgzSNpBNgt/5ROXKX9NSV6AMVDCn4aC5WTpf6sPIaimHgeb
v35wqS853EkDA38XjhUdi2ojog86kcJWBDa5HkVsm2pIYgb8ngT2Ky3qhZ7m5MhVXMsXy5/AKef9
VAL6xx+LeTkqp87Gt64rb25LNCZhk1j1apiZNDKjIMdlNFW3Bbt+dpgNx6hX/EgFlDsSlvtcyG8F
4hLFQY5qx6NJ5M2cxj5cj/JyVpUH+9WeJGBtIIzno/xdB6XyHe6c2dMg8eKe/Fs80WQovq65vdbM
N7grrNajJHBTfUl8yXh0zuyjXJMQ7Q0W6JQhDKgdM4SgXlT9fEck41JfqL6AqnbYOj/l5TQSuuNN
C6P5JsnuA6i5tjICW7AFMDtbav8Taug5OY0qf92szkYkMuvG4MQH1N1C2zp8bFgM+Q/VM5rfjSAs
a7/XpftO1V4ds8i7QgQ7+PONMgNedIcDtFbfQQJV6/WeBKA0P8eZMrDB3V36c0OGNpxvIeTg7rvK
Pbf+gL6cGGwqDi4fFcB/OnhZH+ZA8AYPGDmlTMj12BJbkk0sa8dm8c26ISZ0d3LC+YQHOt5TVaAK
+YJn3be+MMJGkaTvEzf5kLAicO4oPRAP1PmDb+zkWwHGoGiFulK/DUoV1uI8F6ZfhQD+9VtLzM+Y
v0kW9ScokyrdbcEUZS/OZWAIOLbjEsye0Plw5YHv3ZjGjpw3IDbzY5vPWpU/uhnTzojYZ/weEdqO
HGBIOc4MlmRVEN/unSp+fOi+DV/FnZR08k30BGvhXacmBcBcLpsxahct83yvHJRPRa5uMhXpiI8R
QXZoKqwsLhQm5YSpNbN0zViCCHbluWgc91dLpAGmQsBhDskkpPfiBAYnHhnLNdmZV/jk6b6hH6N/
4e+rLI5u9mwtl3CupmK0ZcKWIKLf6c3jtnsG47tdUeLsMS8igYPFWkIWE46eTImH+BYBwuTNgsEm
MPzk6SqaCeNDGGG/oyvB2LFfCceYsGCp60uYsDlbl8eTcyZNtMSOppc7yxVm9gbpZEwIKMz/Xyc9
sKTgqlhmaDpNnwJr/4ttlKjajEgRANQXaqZ18HWAJ0W3KFMDOPuDDSJsPzUbAFTXwitCsJNYH2SG
UNyyNOPgj+3x9+r2RoxQrDV5VUedhzYcYZ58B5HR57o1jmgfidIcad7DTy3KtONJ7sm9M5XvwJN/
4wQKSE9M31mznQmALZo7o55+4gfi1uJWqSz4/NjB3cYHVSgJLWqYCebReh92YtGAqBS+5Fu8uufq
/fRxw2EBIufSple6vxk/Mtuo9upQFUbTrUys64fEGXgpLL24bpr64sUXovPHMPurZ8My8Csgvh6h
5kCTjoKHDbSVG+8nynrHbIYCi87Uc98PusQXdbR81XmDBDNYS27TxHKXEbs65MLJidbW6fHUI/Oh
2sQQsoFQw6JCr/TfagwT/+5dWScUiOJcCNCNKo67guOJw7UZxQhm0hFMzYdVBtRH9JEcjjZp0paq
l/7wULW8Sa2hQVOb9YnRCZ7XSnTA1mrHmrCLgw+Q+yJFa0mVUxA422o04u5bLrR9gufvkJcDRzPR
saDyXGishIiDsb3ceaR2UftnEXP4X5UNayL9xTgTLauRz758Bk5+N4QDxT/aLA+Z6DZQzDuM/C3e
vSTzi09lkPy6fmjkjWpavKtCH/HxbfVEtGHtvPVLEOPDB5lPnNhOSCL+idxCoWBFRimXtQEKR4+C
kt0juTpQZEAArKQRUD1W5ECuCfKCMArq7V+FdozXqF3/1A5ri3gAi4s3ChTJR/Dzh4LJBjWOnEkF
YtXNxEt4gH/gnz6bAHsGeT5VPetmYf49uIgd1n5J0dbmRvfeT0YCW/edIL7ammFM6W4PjfL2sS7e
G8R92hDET8spT4dUlSW5SJYARZnTmjWS/8ewwmiELgbbdEB0r3bVK6Xn7Sm3GB1Y4zCXI5CWOv78
jPMiXZX9yNraE2GF+Gys77r31iM6QgFZcoAOr1Ew5YaT+8NGRhkRghV750FY4/EVVykuP+xF7zpm
1pDw3+xR9ooZXP4HZw4Dgat5890uAGiayHVdL5aQLMjkXhqE0E7GZYLOOj/2R6Iow/hTDCkrh93H
ZttDgJfe5wA1LwVaZSQZL4pLVDEOL9DCrl6yxWLjjKH3lR+wzNXYyRXBSzKMwEqJmn3YnFHJmreU
f375f07M1PAk4JpX/iN8LYSY02kzzRVJkU27HqMi3P9T6yV2BcPxK9ZOrpio4RfpCcLsrpOX+2W8
c0uHwjLOAV48UIUF0Pz2X5pM8FTqMOJ/GzQyZt5XMpYHkHh2SCH2r8cy5TExTZ8mU1ZOXZ6ekOUt
VK9QvYD6stKMhTA1mSKQDetqe5Y/csNzwH7EU7L9i+Gt5eS7B/ymC0vQJd0oSkBWSzcGxsOVZbst
Uh7IPc6lkd34ELzCBf9f4b/whAXuore7pkMx2upZt2BVkGGgYUjZCgIoIqYn4du8jKt306V+5ikB
sDgCjLXDfSWPU7HFViO2zwYkHmaWZb68rurwJEilcwbNaeWnOHdPuLOgEhbrAmdT1eQxcvDUtFW0
loGCsgGJISc55OgqedBmeoJkuekxBLogU0OBm0aErCFohd23T9DJBSprRQu/eVqF/3AGaM4rzcTv
stQQ4BO+/OojJL1uSNaVYQTGRwOmLipdO86wswgeQdZPAicF4j38eUhxudYLy7N1CfzbdIuTyabu
gHk5d9psbgf8Qark5lxw84VSGxxs4rvylJwfjN9XvjuKRdaVCXh1lTMhOoR35j5+lcJZJrf2mKce
zsMAxYqDGhTXT7RfIrcvp2cWNYS/rmAUxiWAsafPSB/uU7qXrzOVbRlGbX5PEfLNj6EqzXlPp6N6
WaBDqEUerY1mqKo3Fd0u3TdWeQU8oC7vFyc/xypVoIvdD2ne52OHxBsfYprHAXqlnZE9a/WnuhLv
Mdx/pWd7wOfrLoMSwmYaH1AYe035gJokheOUUEqxnMb+BeiJBZmwzyVkAx4oD9VqI3k1iZoqXzxd
Vq47OSwHxkaMs8F13VEFloC9PcAAOjvLPh41fJO7/zrZ8E4DhrROeC7YgCMzrw+6FgdR+CxzMQko
om6YXXH942+ITvOJG/70eA4mTL52nS24pd39Ftf367OodJm/+ClBh2ca4w3xK1X1Z96peMsgHdq8
mVNfV6/CnduyUuJF6nnwe2fXGZ6UHx9R565wJyo6EoJ4qX3Tfl/noZIPzy6+VJcIk+3j5HZF8kBL
GXjxvIc2vL1HDyJSTvHpAOEphodwgFqdNdn4BcEt5EJT5ITLP/GIGY9vVEbybUMQ+mKsnEIrEXR5
5NaYgAxxXOphEV5Bird+otSnOU5CzLY7IioYjbKJXUrKLnnAjbYlEeI+PUHlXJekdSf/2Za1aukk
n1WLWgKgLfuaI48Zct8ZXOsHM9m95O7JqOrMTotyA3hnSB58jhGTdKBLRsvWGh0aLADhXSo+ftoK
rlG3OSJU2tQytKm4qMaipD0lLcFxy2+95Vb6FnxDJ7jLqXd26tRlKUnB3Kt7+P1PQrArLTTjYURU
PTgArBsq4x/VBj5O3b6nP/jhhIgGNivJJIgiZEBt0rbwo+/eyijIWD0V5UiWcIaRKxgQTYQp2X2i
k41tPg2E9BzHwm46PVRCcK802bH64pu55SJcwu3A8OMAPWr1FkGucHZMAYBsPpsm/M/UXhdtAfj/
qfb993hO69L+1B1gerPCKE365ontnacg649ROD47QDKyEW2FfDapggln/ALTm2cUg26bfEQnUhUa
xf0MJQXoOVohNGxWk1InRozy5N94MbBmydAI1VWVBKNJt5+FCazgl0jRhkzVF0MqzSpCqBQs0Eqi
7w5UuuSAMBeemFYwjmIDcftoQGe3P1L3s9l26ltTb31MiWNBJ8Vy5iyCBJFAri1Ar8Ju6OpOkYx6
i7v9pG1mHEeKhcrC2kcmf26nyZQwUXoXhSEBnBTFunCapGrLm9dpvaIU7j6MMlSmlw0ryDDS6SyL
5oHH4sgreCbkoMNfv9/G9LByUjqz50Nvf0iGPDmhT1CqABbkixJrraGe5Nj7OJ7aqdC3681LFY4g
NYDc7EAMOZh0IuFLGvIER8uGlySmcL8dIiT/VzH6uvLDIzGTb4dykpV8EUmyk34lWWuHclLEkPrZ
Eg75zbQ7yEcQL0VeWcF8YbWb6dFCkJys7IHfpzH0aHr9UcAY7/9pT3DRjDijN/X03sWJuJtWY0Bf
TpiR3Fx7ThKQGDsjhfWtuJ+adHPsaQJGuqBNiERSrnI5mty9DXRGX0c/2VNeUllEvBSSYJMe+lh/
taYXzH/Sou2fCCB7PTZJ1sa1uQiXfeG8ype2O3YVsoH3Lu9RB2N1/JLvb2Cnmlm7QmYS6fhVqXXg
Z2q+jSK4wScKE7CrNox4fzC2lW6Y8P8QYo/Z+QWlPXYPxGIy/rvaow2bUacBnIQdHXgGPImfAqzP
+eHoF84NzLcKD6KPgJNoWeAhiIKf9wOy6nPdTLDXHhCXo3K5+leAJAD2I/4eDEWdmLEHYdpU1XLZ
NWVvzO0TOKPTpkYoBv3oofU+f0cOvYryLnNUQ4YwZGOziNVofOGDoxyjKuKBweBZ4sR08a1RH119
ZhJvMxALT70fX1YNwVCsVE30blhTCz0U9zDYZHV4pBjXVEFa1j0kQmJvsAhsoyt1Y4ZDOLsT7R/D
T+w4UsES5xS8Uf0m+MGUClZNYlsddZ1clPX23K1S1LLnVsjaCPs2LhmavK9leIm8NVPKMxX5a3kZ
lSxfYY0hBlXCSU7rg1h+qVypVsiHZcBTUn1u5WpXUuVFsdiLK7Nt4yvrsmtMs3qErGsuYF4trD1p
k44JFchl291vYpu/Y/U7aBrHvrJw1mgjk5CT/gA90Dr+jIBeuctjIkEpz8cdLO6cmE3nDomMxF2S
ZfBrLi4jqcbMfaJE0YmE3rKKdisxdz5myFm3PtvynNwtoFJj2ffRLWxj9AFZAWM0CMLUYBOo5/AD
thlM+oxkcuRQhV34GeagoG9FLxSAtQycMXkrX/Mrv0iyofKGL3I7bK+FnS0ITHzjuJ8+Ct4RGZ20
6jvC011zADGcg+CBqWHNSTxKOLGsRLHrnXy5xhdHxo0wS2jkqf5wMKh0c91ck7tXIL6mM63bWsEO
Ob6Ds19LI6CvThSdPdUV+CsurV/t8xTu1HPaZGPXYG8B+ANq17D/YKmcVBCXNP7gUMtTvGX9oDqd
X7RJOs7moDJhvSNXVLMqHN4cYg1gH7njeNansE7Fu43J81EN/BeC+hEexXTHsPdU/9TiBFZGztXa
6ccbjqqFBOR5DT2eHujUkSHyfo6mGJMdJ3KoVeGwdb+zYhIHX4uIKJjsk6C/ZIo4qv0hSVH+QYJA
87EsH+aqf9AjT1dO8jilN65o8otElH3zujuDyJzkWxGo7EnachGi+W4Se3nAOsbvCq40aLHnjSrx
miZZ5ILl49iueKgBFENUZWvcrpJSfuYxEthP5VZLGvZUXLOfaoFnWEh2UeVAKr4NePORXwnb2Tiz
jSNok6fvBe0oBmqT5tpmUoyZ6zUGf9KR0uIxjfceDz1UuOsvKBH+asb8qAyaV/vJcXgsPEwGWzfU
VEVb+3LbJbKPrCt2i1FaAvCyNini5+ro0wxa8pt24Ys+aD1G8SiW2OPGwcBvrpynEcpuYfQtm0D3
ps7uuxiE9dDTV2GW/wHHBIloJYnLbM8t6w2qZhJSAHXumDkSEFgEvi2aQZsCKjeEEQHdHndndtW2
s9ZFA1L8N8+OJliJvQ9cdMfiqO8ehCG+xCr33WX6tZ8eAoEwfToQ5NzIy2iZnwCVqLF83rnmRXQr
dmealAkoFO0xkYfA/I/0WdSUawlzMxqjWceNZ9yeZ3Tj1xBzs4IoKbIAD8vkCT1jszsJX6Wz0M8q
jlw4jAFgd7OyNcJqeaAvz9WAh4EU2wEuE7N8M0ImxYap4Kqk62tYyjqfjN1gWirsBSvYqWMOepg8
hvLLsA78MEiIElhZVkopvTqxj+lFqWOn1a1FMg/foTt70IpAgvi8ongk9V5YVCYbpkEvvPUvrLXG
Dc2pTujvM21RxwdNOzo1faKoawVLZ/s5O6jsxs11bwTkEEAIOjS+WVl8XiedTGr4QmEc394meK+p
/Mq3YVoxf2aZPR+j5GKSvQbqqN4TrwSeYgkDYmA2I/KWZCiQr/VeyXEGj1bJgWCxQ6WhVaKn6LF/
u+31x6T0e7kgs5o+Lj9j90/H00Cf+1w6k9jcgnpxfWTPYw244MfberWraOu5MTIA7KrvE5MT73gm
m/lwXWVwvcCyEdEvflLP2dGq5XqSdIAfI5iYAi8vy5yLcoFqiLWar6gFwZ7nblE8oMQ9iSumFw5r
A0ziR1FrGcGZw0iPbdrnBcS1xSOchsBKzK4IRS8G1W99oTFvEGy2YzJ6ZI+16uvdLq8JdJX0ML9P
cNFpprdNCot/EDs3+xY9JfE5lyNLFNfj0GnC85UVb/OJctZTakF982NGifdOkcedbYUI+SrVCHSp
nJU9HiA8CG1THMfN1nhWiw+plWHCjw6YdENdCRx6Ha2003R339pEKapFh9+P+Z+cBbUi0VV1ifmj
Mt321dfBFY7gtA1vLP2yJsEkx/jWqDmUGbFy1OsgGMW3/Gm1jdRO7goBocZl+YTa6orMfwnbwim7
Cwb2ElyFp7GOYM/90WU4oBvwLS7E95WWFRJkrMJ6+7SX497b5iyYwcv19gTDvN9YsGEZrWLckx4n
iG/CZq5COJgFqwnEPehU6InrVQ3dxk5VFd2tzvdlCQbQcK2uwAjd8M7hSsIwkmyfNBVuqqYv2ll5
Td3Zb4w8c6hJZPUtjTZZnWHT8OFEm4fRsC9xhdP0vYekdLPBhK6It96NdgRSgXAfR9Do0dZk3OJx
M17zYvzhdeYesA5vf2+DQaIwWuD6hMdkQj4Gw4hGuZriPQw55fghvJp2iKFKnCf2nDcp+hDANu61
tYZAKiWX9d57XYcy94NrkQekD9/SdP1fXBBGGtpEbS7QZ8edszEHfPAoMoE2uL4TSL+my7QT+vjM
23zGXuumTC0s8MP+TZL4Ln4vaOIf5Krdsffct8y4F1PV0H85L1As4UfhKt9qbxQM758/f4If1H/z
K9Ws/w8zGqmQtSk3R01+24+10VfbvEyrHbe4vwadAztc4vGb2M1swoVmWvFBfamWZYCBJO/rW5gz
1li4QfaQvx1V4WH05qrxMlWJEsdNBwZyIqhwJXJFM+tczeXkxo0H1yDGjsSM3pGAPumCX0S2Ren/
28G+S5HllJx4NeWxavlFhcm3WF04GzMZgoRpxilicOc0uCLHZncIVKQ3lVLXYPN2SsikDL4bn3fc
MElvSDJCAwD1GucwAy0WAEVRQsKUTJZkdEkNkoqztzZ3KW4R3hoQkqttRikthO2nTt7fapMbQufP
elXi5Q4qm//bx0sFZsLMJzvFisauxi3uWYQH4wZ0jxc+lOU90FXDT92V1CDrOW1XaR7JuKkvEedl
Lwo698Kei/s8YRPhROwGMTvEB4A/szZpV63H1V/vdaNRyWVtyyrJFhYWrRGpfdBDLt6KlzvYadlF
n1cQoujtdA2sNbiNe72mFJMOIBXs1BXX5u/CPVXb8V4mLQMeFVyvtOQ4uQXk0x8vymBqrT11C+MT
REBa7f5E0ql37f2KHlS+49kEVTK+oDBHeK1kzO8ZDeXyAjb/WYR906JMcBgLEqPzhEQoEzwDt8Bo
+1urnjHsRz6f7S1tKm7McDb25aw+K06ruNuqdeN+8WfyOCG6eZ60LGZ6URuPKMYWmWZ+Ulnjkv66
uUKJujxyzIY40RD7S4tFas6vzyQW2ewE/EMfOGKN8wfhU1ybyeUTR1ogMyxZaw8sRgkwscvfD5Th
XUzVtx6mIfffe7+SAiqOiPOUm5Man1GKhOUOqwwWZ9uYCt0TgsY0h1dsKPE60PwbeJgZ7dBfiglQ
n7Ykx8xNlNDKLY7yoYSosFlyCqPAibSgOkSLLMepne5LFlSFkZEfHASAm+pfqdr8/7Itj4MRS5ni
SCU4wlEJKBiB5idjSat5NROLzOLB3kxouGbAgwfS4sI6IY/RIg7jkFt+/gqYnwN1i+fFA59DuO0F
L7diIA7N3ABnG9HcJ5exjraXfRiVyyipG8Obq+UAW4SltfTc9s8Tp+fnTQqY0K81+M5pVQhr4BDM
WHmz1qsGIk4YISmKT+fIM2RZWOiHQxwaTs3euywpbAAvBw9bCEV00drZ0nUuGT56vwGrP1Fy4xoq
hCzpvHSN76Czabww36ldQsGInm1nJQkoy2fOfApr+xuqprqm+b+wavLQ811eeVdxdvs2LDyq///9
klFQZdvR5kQVj+JtH5QR/1TDcJ61ESFm9e9fROloomTpuf/HfNX320TEsjqaI0Bsu4YjaqXhd9Kt
vb8CwnbwYXAN/09k0ub4XZR4H+K9Nia0kRz0gbdt+EDvHpjnNqhj93bDsMkHYzbB+HaGB+JZOO5X
u1/1fQ59gi1V/Y6H/qmC5WDQvJwWjkhJ13IWHARbAAE7pI5P+WTPYTqxgRN5wvkl/llqkkTPFijR
BTMFh0Nsbl5Zv88T8PBWV4eLHr+C/vVTLg/V4yjols3C9U9QT5cQRjLsFTpAzAMSKPvPK2GsciWE
nXQLFFJLYlgJsW1qyyqeJzyo/3ranDghBd4F1obzco9ELqIx7XXV/dKgaeVMw6adKPBXV9A4IO7G
jOvB5VcX2lo2CxNpb1f8lD3yCFY3NCme11+PPUEQKutxVzPGWPnjSyqfkyiiyzb0JafILwg/lbl/
XSfZV77yrp9yF9KWuZ4KMmVaMN0FFZJ+7pmZ0JHD5XztGDZ21+N6zGEFU4CmNNqn7TaDlapz7exh
YRoutEdBO5eBjCix+ELWNP1oYo69MxnoGeFruYlW5vaxlgjKDfFEtMBahcuFe4GDmsJsF7HXxECx
I6SUHAcpv+UwH9y5oRTK8qxJHDn4OhpXX9qyQCtmqulyYZZwlCxfQDJMeuMG04vSdcehLLIHVC9f
eQdz8TpQ1Ik46CUO1Waw/DvGqCBssF3Kw4/wLKjLHiuYJ2OM6Bt8ENy0BQJV1NqziwFHZCV7a1tW
DGry92GwAYDJK+5ydUonhlrrUq0Tf0Q3g2Ffo4PVvaTiD/UMI4O1HYzuvP7XWYUBH7of7dH/AZFl
rVh91KydTuLeWmrYEWtmbIHBiTs3EAt8lKJS7XJt7XOFP6f41PybGCJxsRXZztUMrnul0GOKzPZ1
aQw+/j+koccfDGiN8OKegAFDljI7YVk6/voIht0Al0xHcrdFxag3vD2Vtu/i8Mirq1tYG090mMpE
DeuK6UgLeOsPC4+B68wc5zi8ADQ8m/v0cF6QEoStyvmgsvRo0yyO6gZ/sDqtYwAp6kQZwo7ETffH
hmQUm1WjuAZYmY11uiyYe6ZZMvIUlbmMxysxtQa22PWsHn8pPt3z9CKWUid/vik1oAMpR8jasIij
kPJ1UrjeLlndPGH/Y1kCMqKmgTaMgs8S/49HKWb1KJ3OCxxqvqjkVqPubJivRt7a0p94t4+Nbua2
nsKRM2MTFoccL2zUZ0MbY+g1ekqV33Lyvqn8+XZBMTawsLzSNNJTIGe+1alTPWmEkPkZPg+jSrZn
t1Y1GVcy2p0yXxpQE5H4zTW48VII33BoH7DE3T/0ZoY0/Iu6K7pOyBKtfrJXRRwOdhRmbuo+q2Tz
yI+Ckc2F1rL5UyrkEn16p4bzwsd9pmesOqCAJJGliEmOvf09okMR++v22wF+swoXBElesj3JJfam
35XnRsialbIXDAZX8cNcWwemrDSSfZNa2SAUu9WDg4R+xxcpFmAPVM45UoQuzB8q301pylfo4W/V
c7u1NULvSq60KIyDfTpgumpPFjjKiW0jwPg/quSn+qE8H5wpz8/BZ8XLPGcsbt/ixs6igDIFdIwO
2dOr/yUNGX2wWODYNBYxD8VmDrF5xj5MiEEQ1gsXPyAx55HFXEF8N0/iAMWs6GWIqNbVZ+b9GZZE
iwYXmiLr+cTtvnJXanqxe41mbspI3JCOTMfPldm7Rq7RnLGS8SW204fqkvDt5BTYqMQd4GFSmt5r
rfqPhSERwE/MgfHSRZAHl/J1XymDFX7Qe4XyVomH8nyyed6ABLxk4R2HfISAEuu1ukfjRnTu0u3+
nN11zPgRnSqywJa02Hw1cU+MKJz/xgjnlmaSu19JBfI87PK6X1SM9BMoDZmiYKv1+/He0/ddDGbr
JUnAaMR19HywkhV6WPckkvAZ0KCCf31h8JkkInylqVMXT/PvlICn1jmVHROHAt6zS/RzYuf8NRYw
uyeuuqJyA3bXNKTqRVWHhkgCX2TXIVHLj94dCoMTW5JLZrl95uHQ4JWBkRwnwkGjzTDDohEgqRVo
0erh3xzIVlANAm2irPxbdnh/5PFgP+8qqtgHSJsN0Lw6AV4MkqfGLXQfpCztXd6W6ji0fKul/WGT
voCrYlAAe3geg9O6DfYm/9qLUV+1RfGd0cm7eEGAAVaeb1rKZA/QK7vwaN/0Flv2f+akGR5vEvGj
frX8EAkC8+hLTw5dTJxbRFL3ikndEVfhnQflTBZ1J/1FL1ZHJy5Nup2bdw2+0ktVoV2PLZqRjm3X
YNFB/Y7J7NPoWGcrf38393GIO+XpkxqjU6HMWbkeFzNrHsRV7BA4Izou6QHLV/mIu7fm+fzAZncq
RspWLIO6iy+K4R3yfAp5ZRIBHuLirRfEgppWmIe6W0fP4jS/HNvfg1SUtSpaGjesf8MMgQW8xYDj
GJDXc5IyFl0p5ZMgAtr6YqY3pMr6a8YjSbbT5di0L/n73kHQFIpHzcqV0bkOT0MgdbUUhO/9+to2
PTKyMr3ttPBbHKtuS3/Ev84awKDMlEKnKJhp1rP/BJjVjC34BfmfpRr1Ji1uJ7xRFMV1n79CakNm
Du6jLjHhDG3jxlobRuCL097eE0VUtXdJl0mamr1hHl1iUxGn+OncqPFp3Z1bvBMM5T7AsMzL1em+
WAtavOK+RTYxEI/jtXzFJAiWyAtNW7+XBjkMJmum78/cFAIhKJVart9Zt9WqDSNGVGB+1VcxwCRt
8mAiiMjq3C7AX6/OZoLhjv+lvMJ71AvyNbhn6Br6LWuS6FcPrrrmnf1POJZEavb1ffDgEADj7p9k
ECQ47ZhVXbZuaqrLp2fI9Fy3IJpFVblRsiBDCJGbgL1xoTQalxVpKp/S2Afq6dggHMGrW1Bj9Jol
XKqljK2mjGDXbZ31HY5dv6W50VSOgGbHsrAlbDxa1gXbqhWRavd2YrTav0fQG+t5NwXmg9QKUkuT
BJZxF9ap+0W1bnGqQ3ZU/UZnzgxO34QcG8SMRAFYuv3x3wxJB0B/N8pJi5NrQLBQ20LLZL3p/Uus
Mzd9vliuiST53LGc/YzS4cGfvlOaPqDHvwZ6//nWyfCwGLTi9FGDax/1kVqCl5ldlllAUnzbQW2X
/1yOpxLejZ91nKTcvlPwClMefbzByOTWE7rXeD96icgJd0s2lXVQyek6GxWUGfZmOPgjat/0v+uD
U5XDoJ3b0Dyhlqwb/ED3NXdAO438Z+j1hHZ3VISygmHoTFyzwC7mUGvW2cLxmGTT8oi8mk8bop8O
kdvrz75iipSGWWAYvYjbNQsdK6IxlP/1BblUbfBKjZUSE4dUTGYq4QOnKpoiyeijEN5Vlnz1QpuY
Pyua5ahDEgGT9NEU9zagb/ng49yOR6FIVLFwFsUAOjaFrDiW5U9OYX1KhiHDAunejrqRlX7r+8p6
i6FKnXzwCNFe1h/f0vB4mwwaOomlq2oLrbzODpk0cMljDJtq91kputhcjJuaD4OQJQhM8Aqq9rQ1
AQ2KkQhTvGNHcFUvuLkmu+2ROnqjAM7y0HeykPjT4kv/rnvPWAha0EPZKfxR85pOYbCR9Jj6tzm5
fMV37WZR2QwNc4bg3ktbNZ5SomjUv5mMKFkbv6sizkcJAqnsutTYoIOny2Ze2xUeU9l245RDWvhF
sSuqLEReLUSmkHtAHsfzLRHnubEJOYTp/QPcp+ypT4VwPteJs9zTAp+JG1g8x80MuvNxvKmvkFD+
eg1lHU5mxArVkrsea11KaAOtUABqi9zX5WoETm4a+P+tJwWmM9BV70W27BPX29qEzkdnaSr2Blue
cSl6518NwEb1jDS2Osz58yn4xLlk08qoKTXyxCT92SbUolMj/qpypiXhEunn9PgEJw/qQQ+7ZrUT
kkOJO6HSQOeaui3MR58jC7cUL+S/9fWFctyx5Pnb44XrK8/vx1sDKgU0lLqWbJjadfvRkpADDLNa
G/AKzHS9tIM6TuQ7jGazjoTgz+xVC+Er6/QQaH9wjfc0Q9VGFpG16x4rd/GX7/ynZOHqzhBsgE8F
YWw/BzR5DbPydOsGZLC9zZ1pTYnJNC/Wk+vXC13MoONdke10Vr/1Yy3VsTODfki3sbbY8IBEkaHx
NMJy7O+7u3k+lBpJqUZhjB2gNtXY9yfxTTDlAxUG9NhRVT6eVh+Gh0mRenh7oGnxFRpSsk5hpq6y
w7bjn0QrxeHZyZM+yz00/IhvKDLUh5TKxbf+F7CwxWUzYLkvTes9nm/G50JzqAhPqRrcIPAFIC7o
Nncwc591lfFXW0rGQdAYfYFAavDWa3b/lO+UV49bOHSNE0K9M2KJn9NQSx4gJsW1AWYI/WXwPTfP
R8c9oQkx8v43PHvT0+C1Ogw32yL8lQljhscRxYmMJ5Acb/OmJdoX06v9DcIdLhX1gh+UqIyRLNUr
/xCCM8UMBoxrUo/85bHwdP4h+0rMKtkx3sCfzRQL2IwV09qPsDNlOykInEwRE0M4/EdivPqgjMPD
9lHQM+I0cgWstm6kld6Yug3oEpYw+y8BBwuJqVUHFvHnmSLiofhiEdAlG3pcBCzXeEFow5vHQZEP
8oGZMANrx06DveTDYI0CsTpTtco2RtlOGW9f0qhIA3RrjU5iztdRqLbueAsZSyGGayfrb7cLOs+v
+aFpLoE1GaB2iHHMLRTQ39QbZKL6J9ogEmyE68r+ZOBdCllJtWFCYRkwBhk+OcSKmJ8Loz/y5C3Y
bea5MybhlAVyKGSSvwFFcY881DGUsh50iZARoy3HQtpsTSgvu1KEXeCdcD5Ywq0XV3Q0ngWJMgyl
sY5V33G5qbzGoE2SmNymEE/6XPWMHGIH9+C8jH5rhgL9LE4cix7Z0EUMo9yz/MqM/msmI0DWt1Rx
kG9ycqpDV9ysWIyU5aoKBUm+4iXhzqRJ5CIaMJWX9cBjDqGBOS5x3pRvlcWgn+uBZlzNE1jFmgv1
17BdE4LyoorpnLCnNdllmOVigHq5UcsqMDzh4craUzgLgxyn+dS/EWzQxDj6HaEsjxhVTtbX6sl1
zyeZ5dijjlGF742dJKW7thfvesHzo8eDcc9z5PGcD/xOMVFtC1BsOA9GbJIo7ae/xlKFOp+oVvrV
9Esjwg035Nnz0DHrbyjwRZI7NBoNrDx6mQay1JUN1eqelBuehHEuCR2CqA4qIwbnuuLBfFNhflV2
kPAju4B0knoEyjHlyseSsW4Ko4JcM1NttZaYRLs6lXMGBy8CWecVg7En2jZibLLbWX6NgqwyeDAr
7/LzMKg2iEsDMgR1x7F8qG5gUVfPHUJSKJUYEEjsrmd4/JLEV3v9Rgj4kCwMddQ2AA3V34u1XAUu
LNF3w6zmxcQMKf23SMVzIy38vehDZmiN2N39eNFK/LPUFzTAxf+NW10N+yLjz4mzxgSuFMbAVdlj
qLtYp1mW2Ww7TU1FzwgVInEm703VWzS/rdYKbUdojD6ICo9KLps8Lv0tOAINKOwjAoaMSRBMU1fd
vzL4XIBR+l3i6xLMIf25Rho190H2nvXTgIKD4X4KnEpne6rqVtlnLKA+hMuk1sOcOARcuTXrEv3c
KCh2eyfnESjKUh/rs/APUm6hjvIY+1tmPjFAV+ZWERqZQOL1FgWLrR+ivGEz+L5No5A37stVgWsU
XALWv6wg6eJuYJZ/8Kl8On8nQ8/CiALcfD9wVGppFfOfRd/uyvntuEpNXEWjga2Q69uUMIeF6eXt
u5iQp0RbQJHu0e8XrqcZUOINWBIrCb5SWibyxVox3YxbnlB98cqEnY6mOXSMu9T7+4VE58Slqwy4
q3mo3YlWk5ABqZ+VS86qqPttZnW6AGFrdE41Le5yl7RSHpj07YrKJMU8ImpyY2Yvdj7iAArvUIH7
35RgCDWpFxysUpsbSmyLSeIvQL1ZObJ8hyXY60fTQ/2B6LmEJ0OGvVw4ZCbO5kKRGudGiYz1ke3d
9Wi1HVysTo7r3s+DlLACeB+BxyhOS/T+oW5oOxGUVtJXHurJ30Hmh+0MRLrB8SwiNudWUYMZT+nT
+o1osSCsUSBd2TvpWMinM7V6W1qUahoxLbzfgKCZwwIhFq+aXLXdKC0sBoG3UQdZoUH7VgPvDLbD
FdqpNlBBqEys1v9ClYyMVh4cQB7YTbunh8I3cf4LACgNQq4Zlv+zEE/fXeVYud5rIZmiqjKSVdwI
ObIhw9Ztxwcqh8DC/dvlMrWY0NqgdZzThyYqLC/fuKeX/iMHqIVE50xmss7QvM/tyKaUMQm7byOM
SQjzkDti92nRMX/UtTQYMfWisgSxI+Ht9JWK5iDenQNiiAXEOXsYEKQG7eZt9kKLC50I7doo+p/P
tQ0rqVxXr+2Crk69s2Q45oPlT46REkXK9ASwnDHblQrf3ctKCQMCSthDK20Rr+9dkUGssDBc63/f
Q/07NrsyGg4mW5tWP583V99MqAEZerrPonzZEPra9/Iw0iqIpfH3zJQYr26xvRSi5tD1ZqFZw+3r
TqiXCSLwb3/jnT0NrfBUss329fdUpQSVZY5rW7fmntPxNp/7TkQiFFO7cJcfz02MNVthNqeLFqsQ
sq1hHwfOukyiUi1r5yf5Ux+w8q7UUIVFEL7A7gBGGpejCSpNXCDXq1X8vPh6WJZ/aNMUs+YbfDJZ
9Dr1hTgbN7jEr+XVZ8HwxDgEgBvRjMmB2cFBEg3fxZiZKWmXpH5NCCOq0y1hoTFXqUolc6Ql0JSz
DKlyntGVziN6yVRflhO9uoQqSw7xUaHT/xLw2ZCQYICK8yqKuvC1WbQ6UHh169BpggdRa27+46Gr
LPNhf9XF6EnHk+kyXUJOgIO0mIKWsSDgJQ7iYsH7p/sLZYmTrCtklWcpLD46UbDQ6CyMdoftIgZy
JlaArzQw4eslF1c+NP6qLfrIUUs56IiEneUA7gtzTl0G6CYPR2TOCpo6y6tVKC7kPPsUaEtXF6ZU
/YG9BjOGQay0QdicM2pXHLQdNXwppDP5Slo23TzARs3vXcBMEHUfc3Oj4h2+vb8atzpcBwG+QCJh
2/cBnXf0YWtiv67nCTdrJzHogqUNaxBBU2I2zib5+nxUNI6bnn5pRL34bf/wBr3cfxWvNLtDMT7A
srtS87ZWJW9Wstou3fIp5XS7XMw5CktgxehjTfA9NHBNc6OkLOpOJFGHf87ioIz6TCgYUmQwt63g
fMlQhNjGsNH89irK3kKeHK7b746zIGqB+x5kAD4uDTVlLlQ9PLUB1C1zRYFM8OR1IE4F10yGBO2D
dy0KJ1JqzxjDhy5IFA/h+u3nngyZnQHaGvSbO/KLQx+ToK++nKWlU1gjLGLkpBmH8yG+gXIRDYXv
CIVefgGjUhdad9O5+Gw28yQU/nIHKMsc45jIEcnp2REJCLLshXrW9ej4PfVHAowvYDnKLnLA2wLe
HFuV8vuLxvHXsuWF8E9BPquYBm9iQzhywbFKrUfQp1ITVZdbPmJT8wyKSKq/qJWR/8OnYeyt8O/H
u+vdvslWpSEtQd9uRYPfVnjO1uFMstuTmzOFtQpbVhjiX8pVQYtqzHcAspfhG0NEuUxGNg78syQ7
N+P7tGpCq12btkjet6vjaC1+4/v7DhJvzNBuvqYIsZ1R2JslAgcPGsSA6IlUgyuXob6Tyssn9brn
vkT24qwldMbe1atH55XA/gFWeh6ZGsPXploMnHLD9dURB+mWCpBBZ1hHYblEq9LO7bxqtwNus7iF
Y+kUNluN9LMfmDrNX8UWSUJYmcgsBIXx+So8LX7aqi4DuFoby22eeizxpNnGbsU1ufCQAY0upP7k
QeNTcjPcfeORUtBF587WJwDUMZh3U4ap833uJQM5HdgsezTCm6T9HCj/CfPfxjPh1PEfeGkqZvsv
457Wohgd0yPVvS4ggwrjONtu+jknBsRkrV59zcXmMh/d99Ga5LOU/bCVWZFeRqXxlMBYbR48QIOK
56KK3p1qzhQ1k7+Lr+xtmDIHfL5upkcWW6evawYJcte9ebuQMAAXQZ7y5ihsly8u4/sIz+KI+igm
StZWRCbltWC+GUShrN+qY8ta67x3mGuEATPpsWvl3A6VhKBVEn8noQ4rJV7sWTor8edZ2e5in6Zq
L4TGI/OGDk18B1W7P38vRCso9hu3UWS0pjN+yH9ZpEM7irBxCxAUH7l9dEAe2i1X28dYvQ9XlaQe
QsZAw7dZ75cTVfFCu66u6ODm2d6zsf2guL2lUxH0+eCQzM6EiHuRwbO74LPNI193VtCH6FTA4Pie
XjXgOB2fjwjUjKY8VB/B0VaetfFw4HSiG5A9C2xnPnh0h1qoJLfE4MlbUt3DpULvXvvHknQ0E5yS
O0ock11dPW2F4w+j+hGHTtxK+Njv6iFOT8iIoJ1rFfpRzIuZkKxrszM9TbT9yECAR1guCWbuqEoe
xC34DTVm8g96c8wC51t2XENnn3UlZmLm7UF92+ZLSe+/bKglu51p0okUnRubbkSS26rZ3WnQMB1L
fhFErSlXzB9UKCbCzGAm6EPh+UxzAdIEdZC0XkrbnfSo2OIaf0my6hq5MPKEMDZSDp/WbBXSwcsW
wC5ttZ9HyUTrNKiMbbcqmJxOZ5+VdiHBzHIrlHboGUxzLvUWrGevfgYq80baE/1Mqs1gGdjrbVTB
jdMaeZWv5qAdsJGWANcUbtqxSW7Q5yivxFKHzQQjH7nj2qXa3jqC62ztv0dVz8+FYt746sg1izfK
Z/7IMbfFi8iVoMz6SCjSfNaWOngV9bCvALUcVXTEfPiZgK4cQuuM9u1ql3/cP0GFFVfNzdH3HOr/
kEynHKn2oTe1FK/7HBkAZGejpiwd4X3vDkBu4hxRRsVIDlI6hXZ45lq8PUN1x2iKrGxZNkx2vj2p
U0SNYM72jy81sdZIvlfm4FGK1T7/JP4C9zZcfRlT+GYrpLllq07Devm8ZLd5TABkpVU+Cv2xBcNr
Vhch88MxFGtLkK/wizLSSsl5pQHdi+jsfEf23i9AFwLx9+VVgPRUTyIGEkbeKeHO1oPXK3eolCat
0Q7w9Kn5GTuFMqzKEGOxUalQxl6GRSLZ4PUnyTEeLjcVYmkrUg5dsSCcdJA38HsXOKw5u3o1y2G8
F6CkUY8rjI15hVjzSF/oCdJNwxSMQXgGnrzbyCBC+Ej7OTofUwIKHKPRvMgLux5TwYd1t9Gw+EpA
LfE4757PNATetBw90Mlw2YHaBsyLFQZ/IGYxPhExL8NbTD3QEkGyolYokWzIhTlR86yxBakmp5iM
pxhXPqvq+Q0Hhy/DrS9JE+vcBq4M+A5d1S5ROxWT6F/szrpJEA6G4XEuR5qPs3qJIU2cyQH4tuXS
T5GHHfdHTYXjBJ9x+k+wNw9KsdzvDXmofcpn2+mvb1pXzTDfJZTjitetrG6n83Zj+LNc/dgalql/
mNppSMi7cKWFJgqtrZ4pgpo+045xTF1d39WRqeiG1Ycffoujg1qABAUVhNveM3wcFCKO9ttw+qnb
RCdxlTPvv8PWOP5SS9AAFR/SSYW0GqsDp5wis16OZBERpEDAD28zeTOauTvXi5+zGf65KdOrIzHI
buRYQM2odWVjZltZEJm3EkdJdsp5HXLxAEe7kMYZkGFAlaf8k5WXm5aHx3MDL2dWOVeIfq+PWUzv
hHMSD1F2P0l6veZ6j74i+KnMjhZRcHJIGTQPpGQDNjKmMB7pepD2wU+aWhIUiBoRl/ROxg5Gt3kK
X8yRi1AFkHpCyh/+yi0GfhqHfSHFJbaREgNt5eASMkZ257O1IrRL/Nsm2b+jBuUwji6DK9b0/kco
59NkYzvepciau3IpK6p8F4vhrhNuEjQA41WGbix1JfBHmjEKUCcr+l2LIDZXmirevsikKLo5Cm7D
nmvEF0Er1bZo2pQSTugFWlCwm6a91rvqBKIshczqmWh1OMTZD6IsWEo4klMMqdfioACRFlRS3p8N
50842CujFCRl+8ExZE3UgQtnG1LeNjMwXXy52KeD+EWqsxufnHcg1BU1tFWrAiaHejaKq2nLg+Dm
X9D6O6s5RsrFeJbXcAAwtK9Fi+wTUezN+FF1s+r4PcBvykEn0IjUTnsCBsOJvJWWV6QWVaH3rQ0i
AbfuicBsg0FRmpxJqHgI7AkvDjO4zrU8peFWvkYo/zsIViqjZ+C/3NQSK97vHTnDNMvahaHnvBDC
PwsMCc8uLYhhmSI76vb+xZR8xA2sc+Tuse06CBJI7ywVicMfLJQqcUEt316504D4P56JPvf7vjdw
woqAW6nzlQ5YfEMd6+GL42go5cTrKh3yW5sjxnJXApO/BvzOjAgnEtZmMHGlnKp32BAgY3Tbd11n
iemUrw5EN41Dpry4Q3kbiSNrLZgDTFZjUPsQtfAPR0bBRaJuxrw5qXd8v6AobVQNioDfE6a1Yclg
Rcv6Kwy2RLeqEYNd5SZiP/pIbE9vx2OHwfQJmdpamxWh8XphPA+WeQsqH+1qk/e7f2mPa6NmvRjH
rZ3rQaKDwNtQfoWFdZx29FFwV5E9gbkZaedDY3C1sXPknUeiHNrxE18GBgQ5MNOk9iW/W/5Mwi0K
rVq8NpjnDcZxZjNvwn+a405QscO1jUvvHrv0FMXh8EFPgZXLXWuXMVsdQEP4S0mXn1ijvlTsccIY
Den1MgFKHFCtcjYx3RxCBdUdv7efkBkVRI+5TFFkCx+UgxSFrjkmQW+nOU7cxjjPi21SvnBZbRa8
5Y3+tIMLgZ4agZQPrncmEqKZ9fLDrPYnrels7w5/HRhs9/JZP794TUGSUkwfStCwUnh40+Dzamkp
EmAE+jcE1H68VwXEwwIYzyCwjqw8NaDkyyid2mpvxahe11GF6FZX+vN3GOTKJPGufH3w/gQSX4V1
XDe7HFkUbtJRKyZpDw2FaHVfDYYZZaD59JLBCbp+dY8DbsDCAoUh5mOhG3md8ldbbJ6G66N1KBt6
/xiV2HEgAK+msqjShOrndnhF6pRi/w6rj0Ep2zPm5JF1jWcbFS7Bao0v5WwYpJxs20WeUfSP3WX0
g+6D2080Uz3H/64KA5ctNerxGi8bx6lGE5IgvQ1JFpj3A3M+ViGQE6SfRAu889+JgyI5YE52pjCM
OWthsCt4F8hPBAWVEudMvBiG09o0qJh6Hr0rEAgQ7ljDoZgenUa7oD1gQuvXgl9UYCsychRT0MWK
yzzwFp5yy8NLze2LNroXPxpuyzIXzOTaxXrkkF3FLGZ9M55OSuEL4V23BPi03i5HZgfVOQlCvrYd
BbN80J37pZt+ruCJaXSxeGL0hwGSF3H/RQQZdaTlYNfS+PkqbQKuU4y0Aw5GuYZpoqFlHkdCBj0S
fT2nJu/wYfvHZOzyZHLg4GXEWfZARPnSoLpnKikD5OlH0i8jEx56kC08LQcQ/o3rY9DgYhicfKhH
kX2AWZj6SiZpZH8JWb5j6R9ECWm9qkN0cCwgGkevdZiSQgHpGrQJq2PPnzf5QttLDWgHH+wQDuNT
STG40JUl9ASv2uyhfDmptF7hweoq+JqrWckaqWtVbW2w/6Glh/zDUn9x2A44jT8qf+IuP+RDlmRo
OpSKLkpQBjZLFLtA7cX2hVy/2A1H8UE40oyLQVj1U2HamMZiQAa7y6XGCpzAav8MInnyuFmMzjVS
wOxC6Xakijol6tiWi9YOH7Q+VqdZll+OAu35NZ12zQ0DYuwTigfsHZ7UZVGHMO95of4/F2XkeEfC
Os5qEns6lEN/Glk8eaYtKz58Y50MJgznwXpVIjQmhNRjC/qtR6cUDVldqCsPzJ2i4XlJy+qAO+lK
vvHVTf7oZsKlUGeA2g2crdwmnO8HTxzct5FU3p/ENXJuVpcl8VaaWuECTlYWTbgD915lL92Sj3dd
j7AnkiS+hnLFQSFE8Qk8MhjFwdkxbIc1fOBSpR1OZfFUlSSL6Oia4Kbwamf8F/xtX6NfKW9ZaPNf
slLGvYMTpQsWvAsE2t6PeKT4iECHPNSTzZeM4DBzCyBN+fsoaMGYeIEX6aSmlCHoU5B3QT45p2/F
xaPNxBwRx8qCcbw5vq7J/dmH1cFtwc0yHeU1s//w9a2g8lUFX6hjEL3DUOtFR8DZkgXuA1IC2oPz
oyYA4lpZitFMuUh9dVbp8EEQt+C+cTuaQEycTMbnJ7uJobKc1+T4VvBaPr3FFygvkgZbD6oKZ2es
0wqWHNtPSkyHQe6nTvAQwB8XN1oamMTMz0tMxn59slcED/iMiGaEddQIAktC0nOcz/XGqMzk+oVO
Ie3zSKbSjZgzL7HSdsEWN+oGB9mqkhpsQzWlos6wVnYJdBxNKfNBm9EDLCx79p+NtqeZtP5WzQ8W
YEU0XWIALuVIlZrUDnlNmz9yOrrotHHBeQ5JBVGwG5LIbAFMNcUnYb3QQGbu04P0UxXjz6+Gpr+F
Wwz9rAV0EB3jAWifqdndGFpESqc1tUy4VdSIbe93TL51/BaeaDfIGV/Kk4rGv1YUFFde47QZpZOE
4yEzr5dYl5st18io53c8kGgsQporIkj+upg4K2ApNcT1SIeoWLNbcY/9OvUyPk/PWSRVMFh1B6dx
xBWQrN7pWsdc2sTPLKj3WwzkWa13Nqx/3MdfyIq/D6p8m57LWgjiq65uBo2+MAWeTRUbtT1J8CT+
R7XU3DfGzoOn4jX4I72clIsMfcEcL5O+LChzIdzTxZ/22IE01VSvk+O/MEJa317QG8Uc3zHzv/nN
nbgEAI8AB9Ii700s/PXRd+8pAaAWkerI4l/t7jQB/wxu962VZc7Nv5dw3Gwk304WVb7O2vlQFo9N
Pqv5nVx/dvz7qFXzvImqoqOs8VMJZNXc8Oya/1rmf03tHOydKDVz/KgEPrubj238HlLvrkU17+FF
I6fIGw6r+hDNdbhbUc9fk72YrqeVxXXHPLt/trFSO2aiB18ZRC93KF0R7Z36ETbnblcWe1SI56QG
xsJQUtbuv9UxPrpDL0kA8tCGKxVLyNSCIpbFkuhR6nRrynsgwm0CTd9WBVmyGriJMQVhiodEFGPL
oWWJ1NPd6kqHZpRMjjHgOyylSYFHPJYuf5bixsdKvE9LH6JtMQs5WxhgwRlgLuI4G+9pAv3ptjuf
8qNLiBr/yrTS9LLBexSEZCislmqnUqFiPkxnvZqVSNCtE7sSfrIlDi3+J3vZ45jWGqSIL167y9D3
GIqytvWNu7gr7GJMXk2VWwhqwdQZ+jraMznS2fxG4AIGZ3A/6QO3K0Ua5ZxYGLXJ4Rh5wlP2cfRQ
hzGsA1J6zbsUxbMIdwOsoq8LjFOUXQZGHV+TyzDPM9KcJ5ePZc3hvFNEEEO944IdecV6/+yvXJDs
ujtLPVZy1SR8LPAg5T6pNIJFDvf/6GLrWMkcqOEmY5ItC6K8RIDxePg6OQ5KiWLVF5aSPsnIi2Fc
qV9oue/UDLGXZpW0hiEJO7+pi1sCYAsNK8RfvWtn8NKQtIERRFkc9cwZQ3maXXeC4GcI9pzGzptX
n+UY0hAEX++TkBNqIJz4anRvlroHbEBVmUQNWkuOMVlXtGQGdvRPzNgTJGnz9ec0VbHAno0s7LBi
ZMZc8tSmr6Q597CQGPSG+3K+uKVHnzz80vwIEj+bckA9bLx6bsurfDi203eCE7RMZdMI6sfKoOY4
ibP7mRwTYzLV2us0Q3pwpqPDd52Cvk0YDw87pzcPGHMVZ0aFptLZsSrPF/BxfI04kDsYj7ivGJKz
M03IN7dbwB57uu0TqjQH+Ps/lA34lb4O8G2KYmGiz5JvwFfn9IpZhV9WwnoCcnkBFIlBsfdr9uzn
NnHUozCQGqIWtaB/sSmL4uEnDQNe6a8JnpDM7tw683ORUDrRHm5/IDXZ+NhbXYDqfHKhsPj9iOBa
iG3bv4/wZZvbr0O31CGtqZoK6FS1TenBJp0rFvztqF3E8JZ3nTwhiQCpaqSBFWaL9ODdhwSC+QMK
S6WcGBygWazhHTRFE50sbYhASWmlpLPuDgCtHCbGQdGjfVPG1Cu3gVt/fW6kf8iPM1X3a1CKmvsk
ZOELzXnBGG5/zqBvTzK9dw+QsMTqUL3UHXTvk5GKdwSU70aGSZ4Qn8sSjfbSr3nZRLRJVaAGmAv4
rGbz+dutxrR1etXJHVeWnFP/2lkwJSXrdEo9xzQ7WW4yS2AUwzOvVqEqGmVJQ8UNvZCoZkGBTYCn
CjjqqzZ0ISJunnaO2e4rzCj8Keg28y66MBbxJ4etR4UnMlU+elTQqYBCC2VG2vlOhU246JY8MPcr
EG/nWCIxcuZjAF/fl4Rjj5wweKKzw1aNXyNFBnPF83dOq5zF86a33ZjUg/4OLlqpDWmXhdMEGXm7
9dMvRjZiP1xWx3jQ6IjRd9K9OZRXqtk0CjVSb9qdiTLRA+vAbfWIRo0s7w85z7ih40/gOot1M5Od
NLI7poqIigT3C5PJLJtFBzZ2s99yWluQxxl7YC3ubj1h9vwGQ9RmN0SwI46sTnh/yEBG9kblkT7O
jTImUHLqm4zv0liQ/uzzVpdyhLZBXk8aXRO8H1HbGXWtBC8SbM9DFi9YZzR8YC14Zg4eC/w0dhod
KHBs6oJ2I0dj/DxIzNn5dZXsZ5c9rI27cezg9Br/cc9stnthr0ZO/qKxwRP5MgJ9IuytSaQSpv9o
13QA2Ych4WTLJXr3pxjtbYilc4KJ9LuiD3TJ30QFm+qW3JCHaNhcYsMep2luyTa8MB8haUnvXLNU
bp6Q1uF0dnVc0uk4fS2UjLx0cv/B7tK7fVHYj7h4tbx4Z8PsAgL04/ffS/YaqzmuSwWL4fHDeFuq
FkjLjjYVvRWiCdTPqR/u12wlu+8mzCh88Ud+EOYgiVGhDnh6axb2woznmvuhl/uJMkY4tMiYHY7e
G+dpVh50vFLqTL8LIIUkhPOMf8CRuRCFmQ4MrqhW1wBrHcEGfEwH93e3q3UdPjaJGd3nOBZZ3Ty0
Qn+YmfbVSzzULvhxSSqEuJ6KTaxko9A0V2j8WH+IJ76SzGO00k1/6bbE6saSDLg8WzEK5sjq5rTX
ya194VQ4nRWPRk1rQrPp42vMmhpQSaTqqRUh+8eulhG2oJhInP6wm6P0ZkA54f+XL0FrmeyK2d+u
y+CLvqHo+uTDn7fS+qlbx14lX9twON0g/qgUQP8fzKzyBovoxcEdZ5nhT5UXvxE5LdeattEsSfxr
AR8Fhicr9IY0n2t1JAp1gvYMQSqspS946VU3dAJsx3WNDoAu+m2sSkwpVw/im4+4c8nWtkuU9V1q
U2GEXhmpAbnEVPwEiRP1P/PNiHi6CYkqgqzhy2jUrslUAAod7q8uowvgm07nY2TSsn2t6Bmcy7n6
KPyus8R5K1ln4r9CfAVqIWEFydchvltApzAdXs7GUsZEJqvYDRNuo43Vw10LwE6idDABN6TR0gjU
dpo5LkTVqChIxfTGDhITRYc1nWbPf8Ek+0P7ZJJysrKmDyvPNEI8gC5ZxFILyLPgQyZoS6OIVoRR
Rcuxykp0gLbBbDqxgQIU2FYdfls2vOUYy/H8iiZ2YalKSeEA9akQlk1Rq0/1v2giejhCYsH9P73b
cHUy641cht5dqIYLpw498TMSpuMMauTEYuNKOr8veH4ziWGvVrBNAP80L47vp2vYzyXQ8QcYJ4m7
GjSeqweOyuKoKoWrexS9+5fkaJxFcn42XMAcs6qVilWp8EtN/Nui0qau5wqN6EETfe6sXDXVi5rX
koEL1UqZQw1TCbOcp2UIwgTfjMBnqNHPMscB1KT0f9XUaCmWC3retHrDLFTaMOjOJZ2D7kmmomdb
W15x2y29+I+cKfG2VnxoL6DJEi2zRbXZPE3aHKnvJ1Hcz9BnLt5mMKNE0ckDj3dgiN3w1b/XHslT
etPbIj4sFgWc4+zlTCGaATfHXc9uOoACqZYFEw3QYpVSKcbktDH42jwLDyUuDN2tOmu5UG6w/DqY
O6TayO4IqpPlF0BmZjtIcHKWP8xJ+nfgLcQ2C8w/VUAy8esLt2LeW2/E+P+UPQrS8Eq7eQ7FtRVL
z5OWVbtEUkF2S514S9SjFa2ceYIfYlcVPuHOguCDVg6Bju3OhHRQOfFEb2BYlHLoptWeVER9+hdC
9RUMyNZ0mknWPq+Q7KsSGUZEQVIdZp4/p94uA80hi3L2FsbB6kz7kjxUhH+vJ+Q2qVWNduuONf5Z
5uBhx+M7voe9DTPAYRX9IffCrr7yY1I7kOMOH3etVPzAq2GmwBSX3gU7BH7tj+6k4zojzPdaHrJH
ZOtxuktRc8FZ+6tgC/Brg+Qc7pikqvvtDivvi9s1nIjA6xz14HgDTqvwXpOioG4NPT/rBq0HRzhM
N4m711kTGss/+jkihfcWMHR1torp9Cs0L2+Osv6tqBkm/ok51VpaHQlUuqHnvcZqC+IulkAKDA/h
dXOIR19CTpia+oHHsyRD++cOsIV69y8oG8jnUMAOjikdQRGksqjWBUvulaZEGF9b3ILFO5bAiS1T
WvvQi0+8JYpu8spc8XTJg6j4tW/Id9DmLOeFQ4guFHYkcRCnmhyvMFC+5WL9wAatyPR1NlM0q5je
8ZUMWHum5s+vw3OEVSlrjLzDiSMLWILFQa7XQIThX6S8ByQntdYlwmESEJa+WrMrMCH0BAAeErAg
Wu05zm1+HTssZUDX6xNKm+VOE9aKwn7uIMQfs6W7Xbz97DqXa7jIjyLBFlCvgAbU4mOvL+LDIT79
i6SPIiIQ0WrP+4yo17aLDRc14w8rNuF6C87e/QHSHKn3r1Zj97wUQ/+m0o7PORtV7Lt8I039ODtY
tWkqmPlCMvRWvkjqzOvIFEnjGGjZ4RcJY7CbcTQ4dRzydQJniNIZ2iFVeo/Z6xrmbg0qAoI43GRL
upxqyAC7xzDqsj0Z2+cMhIgnkqk0Yfryi8SbofuTI30elwg6JOFAzXjrmh8kZOXufxUaS/6wTJ/Y
jniK4nCqi8dfAPg+mumRSK5JNeOFDmtPGu/k1kJfPCq75Gj+WI+tXdE6Hk2dwmNn/p0H1g6FW09P
Qwp+FxIKxLyFlRCX292+mL8LIk8Ij7eOZjzT7BQtItdFft815lX8OHU9AMB4Qr1t0p3KYNccmhnM
BNNaLQCrZrKwgNts8PjAUEmckXEbFbZs03x/MkArlyPZOsWziKkO3njTL9y+EvLIgecAkphZPWZ2
3yUuviHv8PnTaZZTRYAKtyg0zsulurI70BriM0dtzDe82pXMiWJab3MBHEEabR+inCguoI0w4I+p
dKRNRQ9DqVx5e3E4u++s4GiEuqArKf0fd7tOqFEx24fC1EL8KOeiVy63Cb5OKM1I9MIJI60RqnrP
zUY3+FWPbckdRS0OL8LCQBf159Hk6T5FmPGyuVgEM+Jnad7NZSfOfS0dS6lSIhbL71gvIWEF6KI3
WE4W+sIU9mOw9NAEddlSqnD8U6riUr47lPBrV/vwYhzr/GyHCLOEl+T/4kQCU/5z1x0lZXzXKuIk
jzKdbpvjGQnCx7yzl/WMb+v1IOEttzGOSWUZ537GaVVYggX4dIAWjDjHHTpdJoHLakh1K5pzLG/e
/J3B+UD7gFQcuQ4BYqqXi/TcA7OW2WX/9z+u4r895iDNIuZGbS7GfA3Ys//1hcSAAsMVkBGJCYke
4VGUHPEpGDIfAhMLjJ0mYabh98z3W8cpLCsI/xZ/pZNU/eRVLIHgFJOkYy4LBMuJ+L/TjdaAQnXp
ba7Jp8yX//KrbwMED0qHrqkzbFCyyLG2ln0xdBsnFAtCsZbTKFv3Uet3X8cPKHr9tS9sQ0pgAcma
9VgmOO7GTcfnkM5CwY5Uhkx7SsspIsEy3JuV40eq6B5rP+bk58pX8nTylZafYW4sJBzeuplSae3M
4rpAXo4106muOEzUHChr5RFPy8Q4Ex6odGHT4ZImOGBS4RhXNZ3kLIeiU6i/lpMPV+AfVYFNtfL8
v5zR93nxuGrUSmEqsWP/hBwWmfh6ttLsvA+MPFYNeCgPK6gmhfwAmRsRdTZZaSOe4gv6DdkBtq8k
KnYI0I6J4pB08QAPIU8qgZytGJG5WORO9t89LTUHtKQnzEy7FVBW6z1UxJ0uCS3BsoV2Vwa1Eyid
SvoXx9goOUW+R7QVcMd9kO0gFh0JH+FoWPDZ2tO6zYDFo0iQOYNc4/rcZ5Qas/FXI3bbJPuorN2J
whZ0cZT7ZH/MtAxoOPi0LFeGzU4ZBn/ixQvdImulFQucee7hORuWOStWPERUCL9yizkLGYNg83qT
nnp207iRbTz7F4yaVWYdUPfojLm0t/O1aascAQCV7Fpg+a22kXnoOTyRPWKM68JICzd/9sFpXuLc
O6Vn/ICqdwOYUSy2DcLflllPHZBYtXj+AO9jtMoGie/TNgUFQd2xc2vcKmwI6Nm2CVqzBpCXiDaW
9z+LiFrbwfzyocv/9a2MjuPhzSyZQgUPZP1OGbtYn7yoy1xqJMCxQO6eGv5S8m8Ve3CAZJHjREPL
mDRK6T/zJQINOpQfZvfV7VWuPx9LfSd3MUFdscry0+YSqE0bSFSZP/sj+e4U+Lv+9Z4G/UMLO7IQ
iFrdNw0bNZsZum4ixiS3a6LQSrkhnAydfL4dxlqaUqDaQDDRQA/rlGCR3OeL7XzXy1ln6qfieXA/
ax1gjqNvqW7FhNwGLlaY0fFTrSpbkLqzgXps4TkqNE29Uzw/M14MwMb1lTAsq75Xfz9enlHKYzn0
EcJA8ALCMHB6/cRL46K/NIqr2NOGM8UZZIbgnv+YG/XjWp/eL6Ly4aag6RZatNPGNmM6Zmlv25zU
Ytu9IZnwtC6znLdwGN8ad6GlR+9K1XJ6JT/bEkXzAeb1B8ZXB+nA/W641z7g0650MNkpMHmNlr+r
/CynYdXL8xlFQXLWyhpFEXk9rgr4oOaluf1jTj/TxOFTGYdKEKzjwlAIYYDzzoL5t//mHRIvIqGj
KTS8f4artSvgO7NFgJkG5IFGKWFsfHIhomOfJYwfp8mDX9514+itbV2i47kVz59lr+YjAMaF75oe
J+n5yYYvKVpSibxFpcBs7Dr1nmESa7URPOCwVaAM5ibf5rlQYlxtICS8MO8SGeS4Ml70A0KkLjfk
IQ+FxKjDGyty9iqswGJDJ1B3y8kP/bEd2Tz0ERHSGuIiRKwtqR5CsD0MSmEuwns9hCqvgljncMK7
BJmd5g6l/AZF6dRujOttuRXSjrkcrvRyXV5QwGv3M8vAVwnsfjl2zeF2W6wccL12a+Euh6+9Frrh
66hJDZI6fiIk2dv9c4mWsKWB6Wj9OeG7Pa5//ibxdeitYzJJlyr5fv5cR0jXjVut6KqPbXF4M/WD
hEjmAekUoI5r2gGJevm+Tz5BqjW4v+5IBB3pDoI4Wqg5weNkRxpp/V3UuJxGZR7831HUQ0eLDVca
jHTNtyO632pRX8bFHo6B96g1X0BIIp1O2HXn392JyvZVbP+6fZN3J8Z0NawRscio0J8z55olYpRy
8yolM/enqzFWiQMWT7AZYLF3S/l0bEnB1OOiitX6hzCgEOnn/fMtb+qxD6cSQUQiXFs5rsM3ybCm
c0Fnp18lrjSl4X+J70YKgrCMIkHOisuiBFr0bwL4datOGUbvc5dAk45jfMt5YpV0F9wupp2Zd+St
AT8WUxOThJGAo9UPhx3z6v0Zp6lZ4iWbq1RGinDMuJSMPAs8oaymdZNymbdToGbhTPEJk+n6NgCE
AcqSul5bpfkpI8psbqHgMY+kq7i+G1oPUdX04dI2imn5+HkFYk1b5Mso7xt+c5v5wiFF/Fazs7pv
JWM25jwg+nEMzF2tKiuK63EjTk3cOREsRGEAItd2LIYqRKKXONsIIFsWqcuYOZFyL/0h10CNOLNd
lUi5t8KDcvxo05uKnuTbRyk3c138C9LqdMAn1OB85hVTTLi9rfop0vWm/dZDYQI+Jn0uIfwHeM4E
DiACnEPAQhTKGl8scoyZxz7qaJR3oePVVI5Fio1MoEO3EnkDnWJy/jwjYf6tFU5YXqWUeQ3Ds9cX
BEVDUe73cTuQyZUdnb/KxUuR4UPn70dw+u59k7LoN0DX2sedJrtDrrY27vlBowH4iLSuKukZXQ1u
KC0s3PlCMzbzOx7X/kT2PwsNSuMj7PRI1pGB6zfSwVJJyw5ArNaJXKN3RpK2otPNHuq2OPK4cRBI
UROx0ClJPY6cI7N4oDQCCu9aPI15A/51yTs73KJOSwwewyxENtB6AXhd+C00w+Zv2OeWMtKMJGAu
AJS1tVVIFbzZNQ+wfRxmUPKrwb2a/oWE43XVpVDhitDIHl4HBfyYfYF3ezO+/POj1BD67CMEA/Bh
+mq3axJZ2mLl3MBEK6Xm0zV6+5ZTRQhgyLtjX8AAShVo1qQ4SXFjb9b+NV0shOnDKAlYPcVoTOXl
aighEvpS4nQnh6Wtur38zO07MomLOdtRTbmGxw7oPyAXmrmA41YtnVVNqnqDpfeT7kM9KPmqRo2v
2VA01yYW/aY4p+tCGlgnQZfF0eEYgF5fpa+6lqryt80xCLor/iCo4DINTnt9cVU6z7xQwOE3vai2
rU8zxCnA91f3gHUSlKQGyuNIvIVJn7Id5QKoa1s5wbnoRZZa3Y5Ovg32cScxFDh59HU50nfqwwL6
ewoowK2DiAtwKOCx/YSnUj7hpIgJKiFHAXbCbXT5ak3QEVIg1g0Rn+VZ09NAe9ZR18D6HaP3H0aF
Y59ZrnDdiNhzj9NC8FT9DK1jC2pPTnE/4LaXawBK0Gje9Mubvud/ZYyluv8nRxr6tmDgWyEMpHYd
DYEBmxVYO0jtPr5xCyd6+PPhlwgM73KMvCeht/RjDOQbTWQEcrskgWREqSG4mqThILHTTJ1b2NPs
n7IzIrOFhuC68oXqitzmN0HwBRo8+4IGw+5g0jgeeC3b37DOMYSpjH4GH4T1lrF48wiISjs3ixRj
d4doOpyV/3Im2feFe0lT5rTTN/vBRgd+lGSACSkltjnTKcrJH78a6PMy85rvPnuioSIrWjn7ZQ2i
jrdSTN+z1YH3cRSoa7dS+Cp6XjbDtMP4/YqXoQZ+KkjefoETXXenWCTLnFEX/uV9MFxlD6oFjAwZ
kRjo4EtiCmXyvU+UW/u0Hwzga/Q+sm2NfXEU5dxljZkv7KEJwvF/wz3vHQ6eV0a4oUMETuxVXPnJ
ql1KP7ConjcAMFjRMlxOrQMjbmCrjpcREPyQ9MFC6MagbbstHkrGts9NjJL3O0Hv4HV4ieIVi83S
YjNXMyOopniocfjC+aAg+tkDpRSDKCfnnyE173IceoTuRcHBclcvHgqg7MMjyAWtH9PYo1Aumx7E
vTvb702zheP1+rKU5GflCpbqyGPnix55KgRXK4PhxknSufw3Wjbib31P4D+E0Gu9uICWXjpx/M4W
9nuWIvoeF36bRzM2sZTAq2l1q2sZmKLXnJJ1G+MW9+sDpdQIOlv7RTtbAp2vuVBvCs6Qmqi0dhcZ
lPts8gIdSch1Rjumnm7W2BwVpywsEidgWJTmLYz4ISAgocyFMClTfeerSTu9uGIfYMnFnB1b+mCC
AM4mBiUQz6ZswyBPGroBS9MQqTqStHGjFy/XQDK9ZIIRHexr2juL3RcYpadYU3NRCAxApEyYbNx/
aaqTbx05d0Pvz5DpS7yHlWZMfYlYSEt7iOHHoQ1YEWVbqmknKXWDFBie0tAKooPhVEyn9Qc/ZNTD
69TQMI4Maz12psHr6y8lBSOWQgQmBoawRVhSNsaxYfMfuXl8Pok08x6dR/mqocQz/0D+PWM/0Dbv
1WkTmyPLezWh3POcaLkeLG0qNTb37b6QG2lFjZVNX/xlo2qffM7B8kkNh+soKJIfDJ95GMzO9ZhX
gxmwOWWhXqjHaVx8sy9n2yTtJi66gdlXw1YKg0YyB8+zvVyribe/6qlf/uvTzaR58oRiqIH6cLJS
teQcy5qTSgDnCHUC4cCCNmMeve+Igf+rtfT4+4UhiZ9Fy0rdJXC1utSMwVRrE3b/SmpKs98eKp1k
mNF0Rr+tYZuOuSIjc7L8v6VpNoFZscuL3kXy6yEL0+pecBU0DcHhqKWan+QGp6L+T8atnLxLLw8J
yw67EhmML2eioZboHMaPgJmW44qHts03XKOGP/QtG3ZUUFUmow3lHpUsySySye2hwCN4vc+t7QxC
VynXe9C7ckml2vf6xRUZgS7NRQgdMCMpkadagXnzCWqkWy669mcA8TqSXS0m/3vqaNrkinDpCiae
eqMLkVgMAeTIp8N7DZqDNh1uSYumQnLe7eFqOp8VVWfzCTrywP32aIdm6qbOzH+CNai+8ZALOj1a
JsoqZ98aVlM6qS6/wK/b+LC9cRUaibDO5mrOCsfaDqqPvot9l+4LTI+FjDOYKH3sBPy9H4wn4rFC
IdfN97+56S7X84DaUhZQ4JRWY0Eda9TEgQx56nVLhcF/XoVaa4+Wi1sd5uy8fVE0eseT2Gp6RUvq
msRpDvxG8VpZY9Yr56KbVWJEG3XW30q5D9mZfz9WrkK0lNLYCWOmd09Gp9kFAd4IA7uABxeYCMGX
d4sJOow5HzPXFXNTvpKUfIaoXFStNKvlwPHT6FqwpMSsEYYaqeSMcDgiUs1RmC39tvujLlQgxC4J
OZ080Z0jQwiUyn332JcDJJHiA/itu8t+QDHABySqg81SlKSYXDS6XHCQfsDgbwdnUIDs9JHfj0Cv
3zKm+d6o8NUq+HoviFKzvD8yLbADx18EDZ5+JZad6X26f2PbOpsMmIiam6m8pShcx5QJNyAvSU6N
+5+eS6+CkraY6DuGD6GRIOZVj9mWdchHo+18w06qjrRx05RxxIh4EaIYrjEZ8Lep/c5gciB7ZhGK
wLt6WDo0RJIBAQTv7j/8T8uhHefRLVQxrfn8dM+dlFXsj10ZhUwkd869vC2cd2AeS2+KflMfoOZk
OVHx387CpAzxc6gA0gLuyfloJJlGHi8vudlf0dBbjdT+OS0pCSug1kEaUZlVe9bYuyZo1CqjxFrC
CZhA+9M4WQXiyho1JwoopXBhegDQ/TNxm+mS/obu6Ku6HgFrZtsgKMgKELSeWXx13ZjjBMlAM575
Joo1dt119OAoVhKlWn2SDYWotItgHn2c4YOmCqdEuleAOAxUFDKusvPAzdjioy66shZPsdYqY4di
WSh9VKd0Phn603S3qMfBLdTZTUp4lmUMtVSFNECeTxZj5SK0CYZJAcOI5q9i98MJBrAOYuT+CX7T
TcxvF0MaLkieFCLnp8qbfm9asQQ7UOjjmcpf46f5Gi+jz4KtlsE9iZmTk9bUTHZKnLPSvIThPHh2
YdtiRERch0FxNDHvrqfJwSqJjtm45xnw0zt7CC695emu/MNjz8ziSDcLN92CxxHAGamPFdR8i0eq
CrIo3M6YxUdM13LVka7uu4VTwQU+pjyWTiKQJABaGlVIwJDPlTPfM9AgqQiKJywczITUej0ludz5
5BglEIzNjahDHb8X03dI/YEMWa7/SL4/rOioJaed3Yy17xRaNuRazr+MG0x4TZrp5xs+Sphjn8tP
4xCwSqtdNMiIvX19eMGELxNj04J720+nddzTkJXGHR9a+HYTQYA9Lpu8fbsrx7dgWI3QeVQStLRS
l8foQYnahtUiMzBMFW17ZgrAsmrGWVRICRDzNWY0m256l3k8lFh+HkbVwciWTYERlNof2Cc3viuo
Cf87wAgNvb396MocrTmO7XOXL3OSxlTGvt6np3S4ScqGht2OEz8T5SXUlb5ZwOMVHTYSsA1FRDsX
mqrOIaX9gOHdLuoQRUnLY2BpxBxaSw7HKG80ssHC/5mK3s4uCc4Meg9ALPhSpQCEVgzAvFvWGCQ2
Sv3NEHVbnAkniGShh9UD+C8JOC96cwuY/Wfm2s8GAUyRHT7JKh17PKykBaG7QsInTd425GSB4Kcx
UUvT64UBemZNZfONBlJPgRuMBdPFrOGW6V7a6fWrBxXULKgRzNiIU7wWrd4Id+m2U7ouyIrVm9mv
KY6M7enAxnqfgwJqZ7nwdGhlmHnOKoGeV9kyvgC5gHIim1mS/EExdxONms8LnatfgqgOCtyMSvmt
9G4EHn77lOW4kHNv8vv2CVIRvHs4nyjVCG4URqZvfpGVecFO2eVbAMh8piKLSijDx5FR2e9QOkI7
dkuPFVR0+7g8QY+TTZc00HxV3QbI7DiRFKgn2utN2OZF4RPSOYtiBiKmDF1de+PLD6fnxpHxKIIi
XaKJ8BwDS3QsPmRcUxqYlnJXxpZeipr2/ew2W8sLbtRImRKNjQsWaNT9yb2qQiKaKHBwJcswHfKh
xjOkVx7XVdj5jkv8VOvcMO/f7ySB4czTtYEJCRyZlMV8cgX08ndUvSJJR5+xl34IBwmK8ZbQoZA9
bXAk9PGWdxCppNZUXOIrlOQDb0PKoc6QFEPUHfnkIOJEYc6c4WVJwFZbUMleqLXfB9gKffrUEouM
zEWoGhPnqgnIHKR8I35riDaUO7/EsFeQ2bu47Rx0MoycjYjLJIdIMO8sz4OeEba0XqC/z5+7WAUe
P2iNbzORMnHzcYsp9JgqjsmIESxDXHhOui6YK5v8nW897wqEL49Qsnpdx1VzPsiMGEzzZtTn55Uu
z8MUBU9p+hodZpYkpfkh2rXTmrjUN6xCDl7nnbDpQS7Up6y/sAaZvckulL1NRp2Ben+69tcTp88d
xrj+vx0nsBXnDZCjs2s1UD9VDN9g2WkwqMRQX6baSlNRKJf/up3HfoVZncIQjslKntpBjiodE1QD
CA5zISDMG40cja3GOx+A+KxDXw1uKMwIcHaTOtWsby4PO2BGe3jKyv6HdwZTufYtLD7cfaDK+L6/
ml2n7cBbucgMddk+J5OE0djj1bhGzvrIqwgrT78WUfGowthGELQaHRReMC6oG33NY7TpQK0HksXK
FCfN8KU1DTlG1QbQPXmt48UaNESdcbgik6Yx0e7CzAA20SM2benHBQIm43pNEgfI72hXS90SSuYM
72um5aSZF2DsAekXAZZNTgxrp2RTHvkN7iSEgaczr0WxXo7rlUSqcmhYOcS7T3CxxWXPmBT/KZCZ
+vkKrQAirbcN+Wc/FevzX7iRZqfPkUiJAUXUxHtcSX8QUGIL7wVo3QU2we7WnCAVmBq1fb73gty6
qsrU0+0KsYX3JaetafI94A53QVXQpCHhjaW9PBZWHVAY/xvJGzIfvgac5fWoiaHxNTfChFvGVxlg
kRtjvL0uIXleIXKVZ+zM8VqAtwf1y6/3u4eL2R8PQxvj3v2L4IgGwbge5FHD7xv75kT4MmQNIi0s
Z8iwlnfGxTVMfKUIa3Tef686SQdUyI05teT6LCZ2F7oBE/Hj/sgcTKYZ+RbTg7xfd+wCCJZXehkm
zIT4q44Gg2JVc8c7i6MNcmpSGgawBr+rkLwSKGDpBCRDxL+fWcCU5dsKk5bgLoT9UqhwpB1UKWOp
JwOHkpfy7/Pw9sYMPLxmPAG9M8U9jUYRLWuc2g/itZovjV1v9akCX75mgB+/h741OhFz1vhRaiLp
aTTbnmcKJ63fMuNroGIsKFt/weqR7a4VSxj+JH5LHi1WM64gGk72L1QjPtPpCAFgBejI8xQe6sTm
89onJfMmV6RuH9rjgd+5z1Tc60X8glxR/SRzbc8pG/+MsUxI5Kf01nl/CG4y8bsBl4ed46h68O39
pBcF1JH3biW4RGrdJNXhpGLPZgoXbZwdTLJN1PUEW8FsziFXOgrlRwfieQxxrZ/SwfwH0Oq86wkB
EmaPvKAuDQ4gzQgYOwO6iVfx6/r0yFcMzTZf03D6m29bZ//QRoFaDOxLD/LoiE12xebSbGNsMimA
frIxWTAqgrHC3mPQ2pRk6akoL+fPDyDZY3dCEwZatRdcmRhIkDF+iEf1lSr5/OesONdDzuWqNnoQ
A5qNZECUPbJkbNT1uP8e0OYitYsaZrAFFA5+G8KGNgrPUn57i7n0m23ewH+t46QqNH83V2qQ8pLi
ZtH8Ndri70/KeGDgEBaSo6ee7p/qcwNRbpGda2B4XthoCQEOYWwZKMKNu/VwnhJe1p/EWPfU70nj
3uTCwFgI4tI+Sc9jZpBknxonmLL2ZjgdKGfjqy/a5j7kcpt+XAW+gvk7QyTWR47WVxI9I0nib13h
lVbP4gipLxRkAlbAy9yME/toceLrty21jKoK7q9PO6RQA6oC1uPqrwQUiQGOXAJBcrTrmVflP2+H
8+CuTZWc9xsQkGymGX21W8zkOatSy1L2nPo9IQ8qLNbHcPpe2ewIP5PQ3UHwhZ78sx/phGIcdc7y
0uP0W4vlRsar+DCz+lUvhAiTIW5EkQkiwKvK0hKC9rldsySD0vuOL8dixucAU6AIv1SRfcqI9NEa
y0CgIxdPm1Wx8c6AhqgzT2r35s77WZepB7JnHWOBoun+iBsa4hohTCmvyJwqOPEJeKCV5Aw1y8Ji
7wdf5LS9gFMDN/z1ZRahB9/JI2vMAnF3cOgWRoHKa9DNzbTeMDCgqfo9QFOMkddu9eP7w25JNsDa
xIORey9V94b1WSxZ9cOOb2vUAfuAmk6JDsYDqJOVROAeBMOoCsrw10O8piJwsrn1vZ9FJgKs4l9B
IN+2wr9SJ/g/atO83n8urrQVrHSLoW1qtRYP1Rnro+z/zIsVadzbvNUUNv6gv/qUk5hemWUDKQ8o
CmUaszMI5cuyvubbWZF109vzetcCF3zgJkdyLmcHO+J43jhuHnj41QeQG2aq5rmrBQyVXPdEQ8E0
STX85Ug/OiL7dqIg/1ajdqm/IIXbnDoURfKKX/zYxUol5ybVSdumErQmBcIWH/fFUM2KS36VZtMy
HnaB0coflnwX32LA0ZQe7RZMgyx5Bz9LwCRRFmHKV4tnhnhxVc1zmW1E82KnMhQl2GkJgUB2Iojv
rf1mdkgJ0dAvMSMhxLHQ2FQOL6g6a5k4r9nJEU+PBV/zjJ5GyTwhaod6sULXapSSQWsMQ+5hmRlM
lwEOlEPnLziaLOBD7Hj2xV+QCjn5TLYWwK2iSeRE43hJlK++hCGjD4bB9TerJI8cIbWKdv8n+xJ8
vl562SDqbw0M0tl7hD9qGal5jkq93HOOzBsybGAbzxYOzlL1UYQrNvaiB0RcX7tzMkg7GTReXsGH
ynWP0jSZ5zYNN40XucJ/E/1GaCGEEi3tULateapr+uLGyKwk9yzZxe7QSzsfg3qbM40/8waHIa0k
WP7ffbmeTUNI8kAoGzsnEw5QEFvr7NulSFWlJHoyXSImUvQC2jOygTaTCi2ss6MyBG8T2osrRe4p
iYVggTp1Z9HJBu/x/Dp0qn4I5l4b2nJNqS+07h5dbieVa1KOB8UQmH6JsNMiVc0dnFb4L6FdF4ze
diyL/V8jGQ/cgu4oFt72DFtv6sr592rbvxP34UTk99QKjPsq+fbmFkWd93qzsLZ/sKSofZjGowGZ
tEYSalz1Wa+HV//8ne9qOSzAu1q67o3az5u9dK+dZ23cWdff3yzotgF9j0XjGXmvlrjD43AsSdCH
dh71Jb6eN+iRvGeOPxrCZ+aqbMqhmQkfmCsracSM9QPqBCyJ3RajzMnPqH48sWks430+MNR68UI+
67TrB06tnZEjbVkBH7VshXr80kueZef6pQ5xhNCxCT3WX88Cwaq/cqxTsz1xj0dmfoueYDSqpNbT
AR/1LmQlyg7VS5OS/V1V/RTwiVfSNFag98pziwtJpH4lwEWYub3ItNA0N0q1T8x0wu7KMfXZ1vLr
I5qIpP8eP+dFMCr84nv9chz0SYZxzJjFZFzW27jDN03AipFiWjVUzRAsdqLg89d8VZUonCRdGQvv
TdnuOGx+OdzBLf7t+fIhEg+j8Wp4q7hCd3b4R8DlVuRW89yNZPzPoRwe0S6g2YODxRsiAmqXzwPA
CO6U/cOqkjht01ZXf3rM3Ps7DPTeveucY6qR0X7q8r4DNrm1lcFCzmoxx2Z58aDuTp0kIGG2oAlh
S6rSgSOzxEWfXVMElYtvZY0ms4ymvDOLgjk9VlDRDNUQhIRIA4Cw07j7aNFxAfxm3Dco1K7vdXr5
SfXj6Sa3bPi4Qfyi3sujB45E7hUKZsLUDJxMXtiW7U+P6Ms706G51sCpUK8FlwCVMklECNz7TGn1
MBd8LAibhdKLcs9fFCRxCrfpX5QjSAI9F+ZccKFJ7IGcnPoQqR0CRB60Z9MV0Gj1HNNLQYzkSu6L
1RUYuK+aY2DqbO5cr/CSfoZjoxTi7k41N5w/X6qr7mJDZpc2Ggro3pESb+NeZX6kJ8bgF7ATjAyP
1Q55rDKK8DYkBP5YzQPynkCzBP103TM3F3Utfo/HxcYzEMohDJaXBxMGWDv+xoJfpScK2MKqd8IF
obr1VsQVPSMC9vkdqUrxD09Urb7hwmglM+xsvHb3rU2nLrdU+40APm+13YRVYuYJI9lrxZiw8V/A
9PiXHV0e+zNvWtSWYKo3XA4EDPbLVMVQy3xsNXSmf3X052K6fteoBzqRMupoHumAdD2s2B7UUii7
N7NI5EFfAF6KM41JJfiCn8xxSSWeXQVLXJ9URJ325pv+ws8po/EtqybLH5Iwd/NR7sfI69QRlp2x
zBRlR6belbFSKqDUn3OMJ7poOcrZkaBQAw/eWCLzGeUSmCTTldCtOQPRPYQjo6LQHImP+uO3mxpq
L2p6SdPJaMfUNn5iJ62Vx43b0djrpSsl5X0SBg+tDTiAd3I7SPAjsP8ScEAmHtcZDipMRg2eFjM1
HkbcQvzarjkxpXrNFmGbG/DMk9Hyyu+jc+A852+f3LMJnjdmVbRH/bsb4owiy3R3yitvcteoNvHw
q/woMIRLpG62I7seO+Z6e7Uh1VQXGfHuPk5zqvV7Cid0JKvC2ZM7kO6X3mADpYtH0tuN35SBqPEO
d767vrGmkg25FRE5h/kmiYRew23b2Bo7vrOTqUoS+eZz45prdKZYWS2Wl4CqUZk0TfTozCaZmBG+
7uu6uhDmKSAQ4XccXTjvb3h+QTR5PAaMYQ4zRtDtwZAFVh9eLZsO9XxdOF+SnT7LCFHdLmhYAnNY
A7APQnkiwrogdpyZN9Pcc88wITpSRqawO3L9oTGbgWU19njy9u0wgAOCuc/zT0s2Yiu4gsY6N5t0
SD7HR2zVWjJ8SoeIINSFgs7k7ImSGFXUGrBn0ZZvJf8/oa9xwnq+uIjxao4am62QOesisLQbyp9N
/lhZee5p2POgZZ74CP8AoKZMT+GRpr4Y7lu6mEKnr8WmyFl6LfZVt5bDFbie9+Kh9I8fpwybe5Zl
WC/YJIAzI7s/aMNZymI9ylqZyTLm/vQGDUr2qZ+QMPPxMb3/+bXATQdnBQD/voha/g7W7IfMIi9O
1pQYsSQC+vYz8GUqsyTdFreXpZuMNkQg8TcYfg6zqqTVBMnUIw81qB7L5hD+ZFUCafgjvlPcdSyO
Iv9Uxc0GtLz77mFUaeKti1WT9Uv3RXZEdVz9ETROe6UbRww86r5yXbS88Ae33CBzS44E2KYytOlv
jOdNezNoOjowa69lxXt5y07egwf5BQvlEh7AKF01dS5J02sH+Qw/v2mU2H9+mghjvZu8a6UOK70a
j0blsrr8r0rvHvfC3kLKR6dvOsIMZFyndtj8U/IoUjx9pg+GnnwVDGZEtyIaOeTcViHsCqnM+i47
oGwa0fLlAyrKn5ScYOuJCUn7M9pVjetLw3HZdysL3xrv1TZS9mdnTqp6AxUjKNIauZL2D8fuubGc
0RE2M10X8TCXJNWRvZx5N1OGWyQfnIO0SP7MwpsPdJkB5kR0HeiaKwuqN9X5QziAd/awTFuzUe82
SUwX+PwwAjzQqyqvGHP97EqerZz5MoVXL8JOVrTDr8WwX0RGvoFDHPDYC5y2WMvcJAi4gNb0wxTX
+Ja5HoVa6Ybxn2umNiTHn2zDuSb9Yca6/hgPMWgTN/FVCRhIpBeHj+hr7XXsiib+sarFlnti16bH
OMwLCTHLUz6AGnHMc142+xn2aJ8FT5OrjADKLmUiJfEbOXysdXnXYCSO5VExCq7KQGetGW45ndPb
B3Szrb9yO2oAqOsG0UTNxOCdwXm7Jtxt8NRiq3YLvilJvv/ZA1wz8adj1Q3JnA3vFbjuwPkuBL8K
DV8BBsCAYnmAKBZ+BDlNZ3Efw8N/eGx4wyIIMboB5I+IvXDYSBAQ8f+4Cg9nPIqi4v5mUKvp/Mu1
Oaz18GdeRwmL77Zd4s/N5fhTTIPh+LAyblPyHYZcb2JqiYr4J9rdPPWRhaK8/Un3IHo6JZjVDV3N
g1YXwd0ZNNpuA6gQA+j4BmXztQPLHG3B9VOZBHvFzKMeH0VkmS4QxQjjgyfhntv1suG9Mlx6FZ9y
PB6Tqt5xylmqcniZ5O23sFVCUEylGzkVO1mjQDkPuJ5IMrakSTOtIoYOvB/c0d7sRgifPj4Pvgul
EcQ2t07d7peoDs7zoX3USvC8+n41RL3e2E9OKxj4PA5YWMiQutxFi/wipW9eLvf/g9TY4DIhNVix
6QJVjlY7M/rEML9bfWJFo0GvH/sfzIK+y3H++qRp4pFiEQ07u76sTccWnKWWg98iOQjKoWcGk0ge
J8+W57KdOsaJD54tPE7rxBSblH5GlgQAohbBKFmpJgCK8Mhq0djKfCHTRRDYUeyQ9I8oJ1dJgOKu
CCrRMEUeVJrwQKrtUiH4U6aAClj2uP9D/1HYsBFCEIxq7KKxbaHWB6qNixtDtm3CeWVDzqxrhPCb
ULBWIynOdBE6eshRFYMoLAFhKZtalgWd9ZfhWoDNB04ingIP+yFbdj8YlmtzkCkVwC14F5ssrhu3
LFlMUjRmBWUOp9RmBkxehTLxDU7hoFXUcy69bs0Y1B4pHbmUyBYCGgtSzfTTT4eV/nVltCHJ080g
eTfYIqcWdeIs7J5ivjX54Ml2XbSXViyaUxOT5PPC4PfdnmemXiwtUqxBTCza2raGGSsVRjn4SJYr
EDuk4nbMCgC4ba2yQujko3SczTv9ParTKZpkswd2cmkSV3bQEqFyvUwPvm6Qb4kbrodTwKzmI8Nu
nytIElFVEwB8Ni/Z9GC/N43OWK8nfKXscAyHR1dO3d1C4G5PSPJZOniMeUprKVcnf2w5AKq4Gvff
DGtx3ihAtJ6+u2u6V7w58yWekLVKPqlv50kfzFRVEy36ab+66sdFnlSL7gCDFOJFSqNbfcT6hWeF
U6+DJRwZ3QB2uIzJIbDnaO0XthvCp36HgblPHDoVvb34VlMoV+saw47GZxkDz7WMXU0SH6g7xe/w
fYw1okV4+kufurN6Dbkm22KKJ5aZww6ewS3UhEc7sl/XDuhCGo0++RbixrgpfZxTV4sJpV1b42Lx
tpe+j+7sOlp0uTgYA/Nr2kAJkWA+G58m92SnW7QGGFU9DIU/eTKgfQk3lgKRI15jxSSbmZMKK58/
ibMHf6VT9oFVgbNuIJn8Z4EzbbUMJzuhABOeW2t+Ox/mtrpaydsw3Abone54/loDdnLT1QTsWft4
hH/BtzTQqzMo6ILPmaNXjgNjmLH7esRHog53LqJeNb2Swjv8Pp64YZqW/XuLtVFPkzNa6gXHkrdu
g3GK2IzWmxlrab7lLtAEIEkJMeSOvEbNrC0Tb0DtQeQuHz2F9xiYnI5C5gFjf9/Ac6nrmoXYkMwJ
01Uhepxhv/qe09fJYa1p9aUMA0P+5baw2tU9GyWFD7mIRP7yBbhsAXz0iYVxfYE1jwz0YzyIUC88
+/XmI3RCUQjuEZJSBROPK83zt1JH+0NybaJKJ+7bmmb8qLKjYeZGL2iSLTLSNqUxhblvewF/6s16
4oBHuABMKHM9eF6mz3LcM6fZPX1byimtZPErFokNaMeMxdAJ9S/FDXv4CZ55DOhiX/keepmmt5XJ
x5siZGy/Zp0dVRDiPMRyXgoKaomhYRFndwpeUtq2gNmniNsdh9klCdhtwM47Exc92Q7Ohul76DMR
iWQZvZ43jXON4gNev6M1o/ii8RA/Goh0GdKTVh47w+FYVluHrPa6yEe0hfwtHZFey+x8XZZvaBfc
yFvhc8K/yKZGyh8LQRmG11k6sWhhjHhJMG02o7LqBj6v1llb51sbkNVXI5khutLLiHFMiZddk3+b
cp7yck8v0tvf40DI3ND1e4zYUJjmOWU3uh+KyoZZppa8x06+m8CJ8NGdsEuRfpgIsgCUFKQhaQyd
xbkFny331cjrtr4SS9KvWY2/XrNd1SAaIAuhCF6CTRYWCmaOBfEYgzARjNTkJZgrS1eZY5mPz3RD
lPvKRk01h/mUv9OWGz9KWSvT+6ZPzzKAz2vOKjmV74RWwDV8bWlH0CxAOYhnDVjli40HThP2ZFlB
i7OTE5kHx+qwbNFw1FbQ9dCSLmxr14f8h4qhtFsJiqjpthUVrPs2Na9dNxvAyyP964GralWQnkZK
Bt9d32UY557wUQ3RRjJ8fbeipw6E0ZZrcMuBf5GJB7yx/q4mLVqEyn7SCjK5xgzyO+dUZpqO656T
qgPEubZVL9nkEgvHTuD/b5bIaX2iZgZ98NSwf8evUDKoDStEh6ZGfhNElAPf+g83nGjP9RnWvZ+w
/OVAbCv+ZTANqSGuoR9XTRSrbV5vaAKXGlrS3P+dfggGCa55ka9guCGPNnJWt9D86i6Q2Y98fb8o
hNSVJeTfnFDm8xX+ot1e1hdazIg/cicpFrQO/84u7xQTWqhNtdgXSkV+FL9i8L3mkby3Y/oTGlWv
0ES7FNqL7dS23AvuMPy+ZcU0J+jb54Gp2OAvZw+gmHuVOt+4tH9sCO/HZTUEzAEFVVKUcnRoaXua
7xZsjZPslQM+JPyt+k+DejtaMVvewpNOCyZuPxy3fEL4emeWEfV4EHxZ9IcdptuOdxCdOuzrs7ih
+7VLou0IpFAIVvHA18xhyKu/s5BPPuFXdvSBGe1GJV7h1549PCfUJDOGQAdqAVKxdrLZ7hx/7MEV
GtyCNWm3HcC6MJjDENa4fKMW+tpiYZyeor/1CoP2Jfh4ye72SsRvEVyTg4TMmJpZE2vfSsAwACSU
kuw5czNYgoHnqMeOc1lm1uthn2PiHuiR2j+mLuwmStNIBqa7q0CTUZSH1CFK+YXgJFPTA4rR/omi
LLV2Y/Qy57O4qUv4QCtBQTdZI9eTYO3hx3ijQFkhmek3MKBuSjOyH9T+wyGU3pOdayKF/ZDpx6us
lf9UWSX79jSU4N80FkBy42tenb0YZVbMf2Iwlic/RoD+CSz1K7y8SJC7azzfAvnf6WE+P2JB+KPc
zs13sQ0PLkB11HtwGCGeFQ5e2auPWDHiQAFAGkHGoLb5WtZE8EyU84VwZ+fUUbL2zGlR4rXfUEgv
tVm1CfSVTpTk7naEf3EWCPcJyGdvsF+G66NAxS/wsJToB2vVzwZVOOtchrTyn3PHXLpurInkrhKt
o9amaUcSOzYYhIEzNsmdzJNRHABjK5lw7/c/k0SxhTrC7F0SH+tiGrLKPqLiUQtqgjE/DUm2QGrx
ATS5KYT/jfTB+EoAQran5tNLpqoTElVnoJOgNib01dSN73BcbUZPk4mmYH0fYrQaBaVk64eRNK7R
OBjwp1Zb6XVICkJsdD1/Y6PZQhVSy5O5V2PaXq46LHTIpkJw4S0SsVUKT1Vgb7WG7STuxRdmf4Ls
uM7j/evLOVrou7Sa6xtyMVBEi1lm5WShY7ZEB6O+1ZhNs5rpV3IWNp87qhGnPGJopRIH6OXNZyJ+
HmbK64xag3tHAVHXQvV9oYjz2YL8v5XEywajKQOlzrrb2334AwTQSh0y3Z+zB3QbM5XYcW/bXbTt
CGFNakDsfAkUBQAb5ffuQ2th2eWcgezk8NeTMVT0ZkUnLXMCQs1UUSBNV6ySIrvZ0KQuf8yR8ZYT
gW6BnyECznMXvpqP22Ec6rpkMMGUtREX4Uurn10rZkhCIhNYSYqoPYhsxHUszCf9HaBsSft7H67/
ia+xqk4Tvab2Lg7xHLqtjYqdI4Dd8gxzzTGhGVjyXulUuDt/BYc1NzV8h6atZMFVHdt8FKq9OSz+
h6x8e3TAUf+PQxp/PalYO6Ih1tI+Uzp2qS+jHUq0r+acjQj0aMO9TMhVOBVHZcWGDLApRSYJd/vK
5RBQj8uQ4ZiAoIwCoPDPQ9LWauzAb6WYtJcj8/52uJLAHFbY6fdGaCtTKp/XS+SBWjtL2gLLT92E
cLSk/sbtUY4g6zL6nX/93acb1IYy5h85/8sr7kmcWcDmufqD0QEoa1P3SyWsyZlqFJ4BmytgkMD0
5nG9RDBoL/ENebm4f/Ks8SrOtIsMOC26TDBQ07TUGPyUjlm7/mvydG0XeTMD155CmV8MP+3t0uqh
Wg6OSPz5sT1UguFmPStOr1qIwGHo9NmYy0S/JF6mocHwr8e4jAKwuAzww8zLiGbN5BZfFjNJtx/7
UeRsK6KyC6NwF5qdSj1IZJ4/QQWn5VDgftkUlIhtrYoU5pE1KUU/KFCEE3jEREv9SxCcaPq2Lsjz
Sv4Jk5lUnPnkQaKjec8cIqAoqR9rrt6duPEJH5SK+7M8pnk9ERplQ6/6+sSsumKzNl+qrAWCcYqn
PnEyOTtzG9gSBfSnnHd41wEMeX6NIV53aHATE6g1hHP+nyGNOzsmUBFFSDj33Mtc1WpbZxf8DE4+
DSKfwifZ4b+AGA7jz8uT6pWFliIyU/lMPXkxRO5IR7v/msmXtEWRgyTesnRspKjfErfq0uuvYZis
hyuxbsc/8MWqLMsrLy1Pfioe1xoB6ljtpOYKhX5YoWJWI1/9ioBiwvCJHq1ii1Ry271pciZdYQN4
8X40bOlmTLeZRpVqNfYeEzaMLSZ9E8+NkmwzY8wAx3eswRMSbh+5E3v0GZo7Q2GJlM6Hjtjz85Nc
rErI/5mfyaDBhLe4DW30x2i6hTMVcTZ7GX3KZWQKVdGQmBPzVD51mtdWIsBkFTkAfrI5PSFlUGUI
tAe/1p5MMoWYK5QJzpevOQm8jIwGu3obqicLW3U2xWGAP0YX+JGtVwaRbo28OjLuLJcTrUjzGQx9
4/JQl2MdJyQSVIn9MYDf1XayfpstGHv+JFGRjulghRF5PV2ZrajumeMop44NrtwGVgOg7loQNE+C
/mUOqzDm8Nzlwbc9D4DxOAYqmcGT+lp8gxhCti3DntVr1X20ciFgiTZ3iT8EMy2FwgGUPflAGeYz
L+60DQhv+RZQgHG9FawDYcNDg4PY6A6ov6tOyyV3HTPQqwkJ+SnoNyh99bYKUR1+vGgsdiaHUdgU
u47SGA/KGmKj5r+S7V0F9+iuBDIsD9tHsWJth4hsSUH9Bns77qHakI7O+O452+F/X9mZ0tVzBjzy
pEKu2CQW6zb4LEdCrOipMENLuC/9YnFOQeO7RzdfuJchnK84wiTYTIraDPtZB0EuUoJiOrTRSKYr
0HoKkNEVtskTW3q39T93FLCz/4ooj82SK29JmclbVk+5ZaCFlhSmPdCodHY2Tq2kyAcCmtSgmyIz
/N5kSeMytYDHnOkWr8hfAk0cXYs7H5kVrC1xJIsv0ri+lHzWRQ+N1I/0OyjVKEKEMu/lbHCII7qq
gl8DiLNWp6+Xb594CnoOleRxf4yepIb7hrnGZDz/QNuQkCGOp05M6xZcKRZiNE3noPi1Nq4G5hSt
9+HsK2Dv7U28hiEdAXcDpXC+U1sQHw4zyybsWxDTE5fkLUGo25dD3Py8nnmpnA+C75HFFIDj45sH
e4zgg1OmixcRa8M4DgJicz0bZ3NOLdoOkpeNgeXEXTfb3F5R8gJ9oHJdv9KUuWEsPoJPN1skgm7Y
FIFpfjtZlPscTKZD73wbffpxjFCiSFPyzHlF2J3UvDiML4svAs5lZLyl4tc24RrQFN/6OjRnF1Zr
wWXSb4o/E8E4DGozFogIOq2wX88+bRPhlsHs3lhLu1trCB/GWENncyvvqih3JdOFoonoza1PBkUQ
Lu6UL1gfQpzw5IeJ7Sz3NcnFPPJbTEtRKXWLLyrjfnYzxzXV9yjdZBhMMcOYnFcWQaTza+Uja8M/
9Wvulbr3o6zwo9NRpMwyqoTnlc6LUIGXaLZM3mpEPIYGLRa9zFanjyJIQAKNkvqFJ18dtV5GwrOV
bb9emmXBOgcY589syEzM606K3Hi3mmdF/Y4dldoXpsPCOhOxi4HpivVMYl9nz/InIk/ImrBk5cNB
nJ+cetqk4c4bZpAgwQIHjXEFRa7Y//q7CX7yL6lbw0A0VBNgwbwS6wPKrvivCLDM7mvzDGUA48eB
BjtyDAWrtj7/hVFqWgq7pj5GBEkRg6BIKWGJsvhVx3+S+Et7EE2AoopGGr1eRwOnud9IX77MMNDB
8PvrFwBrfapwgHpH/KiiryqzqlmoQirVBVxJABxr94UqOa3i6jj1fBazQNzQi58Zvn3YyhhOBgL+
Evh9CrMKn9AkW15JqCYzmo1Q5frdWw9O2MLYAWrtu7x6gtwXuBnAQzeO0vgcVE2mg7ctY0K5PyrI
AAR29PYYCcwShwlEDhXX5lSdEgbDce1+Ah9n28Y1pb7HWRpjCr5TQ5PlEzjMdIMnm5KSSH3AkGF1
qx7KmrxghSIOR3IM+mgVbgHs/NkYU9u1EV9vo9Ap4qYCoXzXC0qMbL4CKonR6qEJ9GkPpfSsGWQ2
JdIfDpzwPH27IHiUj9UVqRNl1H1jca24o/BGnHmVpKIDfp6rZduQ5hZjnyGowQfzhJzEMKvC2l0Q
ZLAtbwrXhP57pO9NQXT6ns3ObSOO5zR+LTnVNh9IARgNd4Aq/C5WX+/CZF7OxTohLoOInfxdMe58
IhoR6SWI0a/33L7bYqM6ZLoLez7NVhuoJJrq7l7v8fntOhDUe6qWvd+l5pFY9IhyQEilwEsRw5rC
/EBeBcdFk4ZYDhFAooWb2ysITGDnZIZjQOdSXuAwTcpB+7pMKWaq8qhFcvsnFWyT1bdRMiNak+x+
yiKDLnLSzz+Usf7bTaZDjIPDKoZng977MbfbNyI2xxNXo8kmpj+viK3HiyoZGyIUChvD5C0s9LvY
Its2xDDUnZw3ojFK2EHdOubihYX5mlHx9F4eYRywFV1J+37c31nrEHx8fWzltlZzpFtt7XhmrFgI
ukPKCEmAKmLhWTetyy/4fdCJZFqoKJ2/hAdQLGALS+lmcGiX2mvpxBcM2b1ZAx+A9IT3lBBkuszV
OgcPW2r//IUPRqIUgZqPh3laf1ftqh4t5inY+of3X8J8UwjQC8FjlcujL5b3i63DLQO2JuzvN3H6
8N7+ysNQg5Cy3C7BJAg51rEEY+yzuGv057gSOFJ1Wsc+4EkoRJwHq5EFUiv2s3TR0zPcQRw/+8Zr
1+fG2LOZJ37LNZ1bvXNe2ytyUl6d5Hrk1BZZI9s87lnW1socJAOsuRjrXL/NEoE5UHe2NoO9aWZ5
rSWI0wKZmVTKXeSzlKXdnygV+YWqys0bZO72Xz+bfnb7pD82By7Ko7Ejnors3VhXfj4zfyhNF0Hz
o/LITfczi7R3UESWsxk0NCjlgsmezkQyMuNlrSi81Ww7slhI3GE8ItTm8ipY46A5alL2B+PcMqAs
8InxYw/JSmCRCW/WxopCM1tvc38TQ2TWWZHMlIuR+PmuzHG+Cg+gObVS49r2XkkyOdHyNPh7moT9
IsxTiDeLSkkfcORPKYRVR1KWnkZiUYjWW/Bxhxemuopqp8Rg5hU67CVQ0KAUGdvpzfrY3CJjzz8M
T9Nh2LrhoccKmNGtE5syDLPPBW2Pwr5oV/GhxNFCJlXR7IQ03aETlhoip+0mOGvsgai7NPVd7Unu
0FKc+dGBH6615OmQqgw2in3W2X4P1FYoib1DjfasaFBWmVEwEbigAIDIVzKSze0Hw++tV8z6qsHg
pajXYU91xtJiDQU7B3xoejaoTverQ7UQiPwmw5D7l8tfCmc3+pe3A4B1+Lh5S7hzdL1KRNv4vCxG
KfWOhavwmwXnnUi6qZLYghZ9lzQl81C9tXetWkLqxXxteudV2SW3N9QPqb5o7blCVhxO9Gqrrj5k
Nm0zlWRd2NmWZ6tOvZlyEV0NexTS4RfqvzeMRNxzC9EH0UTcHOtQozhZEkggI5JwLhwX/LaJdftH
Y8xGsocw0aYC2SsQ4JF4++JKtFKiSrCgQE7AU3l8/fElRrTJVF1RPIP04zpV9tLb13XrmXOSKRt6
ZiXiKlqa+9BlpRKMwbREjrxUS/QWNfx97uzpHedcTpX8SoODCGRRgmd/zwhYLbjfPktj3ISVeDeS
gQJyccVsFi3XB3x8ol+tmYE9l4j609Rwc4ux5DBPYS0jAOAySG0Wh5pucSBc87gJ2qGV7/l3F4fp
1NVg/i/98V4e7/4G+NLhkFGyaIuaFVoTLR3SoZg9TCkZaZHOLDPahD+ph6bPKVFFi+Y7z/ud9xL5
xJ5ozYGQfxEdwD5KCTAB3ndjMO58fHVYEOJbnVERJxFfIWJT6G5VYIbG/GJBJ48MaJdQEQkuk7j1
Rxk09jpyFK49zhkGm3ElL2hizEpY5X2+zvxVXMC0aoUila8mmHZa+4f5mn88U96l81scTgyKV/DL
B1pxxWMEnEdqVxPqHZhD03PLx4pGtMyHtShA1ua5gERKrGKoxB5LN4rESvRxwMwZCksgXxFoLl69
n8lmXsCv7DH9G4PZYXYw7rtmj4mqMzML5JqfZI1m3lXoc75NuN7rgmHhYsk3PaeTrrsXGYlGstQn
bShULjGGA7zNC9TclKANETJoDejubVuWfnekukR9OyoDkrFVe+TwzADaEKtmfzgLBZ1OgQ4/LrbM
6tOYaWeILAQ8wDatqMXikyv/UrU9gBhcutMq0ODStNK/6C0nLdjuRXiTtQETYdkYw7RPNmV3sVur
Q/jAHRUGFkNsdiOhPks9bcgMSn4V5uF74b+Zs52fmczg5Bmpw9PVPjtiD7fsNJ0eoE69uaBhXOi/
cJhnT9AWLRaQQWb8S871wQE6Rd8nCxt1IKRe6k3T7li2HH+LcBmRrWk8YXmHZA87Ou2NbCEyge8s
3jGDQsZ1WLgHs/h6oNO/OjyAsQarVUBbNHscL5mdxP6X9bFnduriAa21r69dNuN2Flk/XntRkxdL
yvfxhYG1ZdBUpjTxihL2yJ78+ealOMJdXBAS8pp5obW39xu3sw9qcHHtAlwNtnQN9EI8cL/pnNGS
wX6bzMSu7u/83H2fM8c/gM+tQy0eRFugqO/cdBJ/m/atuCwIb/ofRpY3FEnbCl0Jxcaqis1rWzMU
m5WXd0x9sjN5+lVIgK5e08/VgJdtkL78KPQPgO915oD6dbAb2jvFSHiFxQpwdOdtjwc1dF28FcUT
c7CLnOwYWm1NjSggHfwse1D3z5PWYhQa/UtTVb1Fhq16RWzjidsKbfvxoDvYPoDJyCuBZFRPEGm0
TMp1O2sppxTKRFOBbFpEnr7wiHTkjxAbgQu8kZGV25GTJf4VkL8YnEVNSWo4Fr1Ml7SieXxMNzkW
UlrMc6Sq92a2t8BTGZ6Wh0YjUJsCj6q0qeXAoitN/NAe/kjik73Zgl/IQpPIbBvdtAYONqRWjdBt
lyEXlWd1ZEy226vn3SoZhtbBgq7oFR8CS+8mduWzjC9GOsODEUgm2/N1oNAE1tZv1LOtIgvdUeTw
M8bvO3q0WbRszDAs4pbYL0nKBA6qsyu3Pl/CKKxoJDuCOlBA3fZlGf9Ai5ioIsaNb7nj1S/sj86w
99eCVF8uxGMV2vPBULfITHDvdy6S1V/I/uGtFc1I7hzwKMRc8PeI4vjPUHzWdG2gSEvkdMZQbiSG
CBmFMYApNpzx/d0Dl7HI8ocKF4m8NCvJE3SFV69SNl+UxI8JLVv0VmU0P3C+VqIcbqEfUB51Xuo6
JjMbzRKY0UHTOl4YXVkqKegnLD8MGBeKZbqfzqkKSjRG6cR5agXdXdI0+nHZ+78hXLrfbzSldcrY
EaMKPFzd2jWvL05c7oCUCUKh5UcWwQWAayArfF/7JbrSWtzQ56nGnmCwRo8Pq+nCUJNo/P9t5TZx
ZeY/aqVGjs9XGHnPNBINWHhNfFvITMFfWIRVmMoLOlzJch983YoDLdBiJGgJVDgUqfGzeT1rgoVi
Es7PuKIwlVBodhwcalNrZO1nX+nZTHuXwc/G7I8yKuCRe1sD1CfevXMd5Udx/c1nnEYovQdltB5O
qc37J85k4fzTnsWCNpvdUpE+bwsMhAhK5PLLVWk4dUBAladu5M+n7+4dBMNuNd/crtlIGpn0IoFH
F4mNbiDd8altlN/TWR0uaN0mQvkNuyFXKcDHddFjslyN5IdKRmVo1jRwif/PjOUDkpKvoGupdYCf
ZYqjU8UY06E8ZFumjxuvVAhpWZHGr5jGndz6Z1v2+b/EQiIYVk2m+L3p1ehN7AV+pAZGjW4pf7SK
BWJRWhPFUoxlqd1EY6NA8SAJwZkBGHhmCkaQ7z+GoYfWHPsmAtP7oo1/P6wWnEv8+2phqnbTO+vS
ipiEvcdPfx3BpPQlb7MrOpwybxlajTqMEUCcaQvrtbW+z1DuRQ8b6ohn8SAHfp3KyF4a1HdjPSVh
RbPHFFGuGi4Lm3yZCs0towIw29fownDwEv9CPTfHGUosOpjA3LC+Pc/1L5muUsTBjQhgjDIgAQD6
XB6ZaGHHBqS1ICtC66nzRh8PQL8RhhT6zSRA5F1relOMtuTAKwq4OwevTC9Sm8X+rMZZolSVzdR+
8M7uRcnsk5epS0xgLqTKdteuX/jUQPzYpEB+4npC3Y9sDbnr//2vvJtVV3pMN48NlxH3lW5/9+g4
omitB7lpFEneQYv+L7UUZbK37avizPTEG1F1dwi6ZTtjmDE64O2ypF/2xXKi80TBtcj+R4yoMWPZ
0KsYHy1kCZkHhYE3qAb5mOjg5ZYfdd274EYFV3BYxAt1FnsH+qaG4OZdcu0onvtU091xneufhxiQ
1j3wumyPfe5ugAHzdwvvVfmsZKSVK5F3E/GcTzH0S0foFbjIqBWcng3ANL4eS/oy6fzXQXERVqme
5IN9rwZkJmQqoia6cxmVzDc/GdBdy9O4W93TXtCU0x+LdIkKCork4vhViMtykgkTx4qnHTQCKTh1
yN6H+9V/toEWeOiMaFHiJJ1cmaXTT66ZFc66/BBU9uMmyryELkhfgBsSYuD4YS6zyLf+6bxmohOh
CugzJ3Ryu2zLMHg1C5L2L7IJAaB0Q9OfK1ajbWOF9JvxCZcQNwRmJs1L3dV59G6/r+vjn4p2l34j
OA2slj5g/gSeUhVcaobx9tt2bdq0dDPnuElpZgNq6y3NXhkxGc2AEwPckyfWP0hae7yn3wOTyn+H
yK+sj42E0HVUDyuZr+S3JPasdcm7OXhB2OU7JNqjAxLtKJLLp+qjJd1g7+YkLzL69kIR/BEYQNn2
iD466s0VcNeTUYyZlYWqJYC1AzZLeFoQzX/7qvUhxc47a2cZAsf/Hef0asnnYwiw3UxoxLsVmfMi
lOxI2Y8xUkzj0bLl4Ro8yBvhXhJzrB1nyEVph+vL1mz4EwsbReDZMzWm3e/rTiJG3zmIyKlyLO4q
/pAm6tzqER4qJNc6uJbqI8UN3va02jiB2V2JwYEPD//jsQcdndNPULZjzNRAEgOzPxe2wD27VY0+
mqhQtAf+09KLfqIV5NsI/2gW6gyGJ9lxwB1f6IoVfPMG5ezYeVq3uGoj46FNhmTtwFS4Y+f2c+SV
pm3RLLYrH/evftd3G2IVMH2UbFOCbjmBgYXYZKJcbkCv5XMzcWhSqw3OJtWCTbXVYfFkx1d66Iik
DekxQ5Yeg7LT4Nv1QP/zX6gsBKvYK8KOGKSzwAU2ZQWN+ZNZ4TOvwK+vBzsvG42ySvoTqZpkKqKA
ffSssM+PHH9akmdn8FjjsxdFRhFUhJYmRmcqCqRiABDZt3asIEuR5zPxrfSl7CENM5Bnc1wh9iaU
kXBvMRBfdCCJjc7v6jZwaAoHIc4cYJkP1QEeXHVOCsBL/x9AfdK2PxvZB04btqgnAXIATnQYNFK7
MYFVsLW/P9cDFq66C6E7+2v4bu9orK0azHCxaYJdWUl9RancLkYyza+dsRJWs19a++WdpJ9l/Seu
wgpb8oNJ9iO03ulpHbNaOwhcQ3h4dwOybWgmHAoxhk26I4n5RWNIjlcZ1jsOZxEsd7O0/Ioclm0q
rmpqcJTDAdj7v353jNF/n67YZDSVuNiUZIzqkYbUgzHrrdCixueOTM7dW8h4nm38TR/7DvjTe9Es
mQ1nRFcUf+bGXoXG9/m5G4HmBQAe7EZ/jfV3bj8c+Txy00RBpN48CHS/a2pVYE5/KLzCqhWodyv2
UvuwLktsiDBElVltDXUWqXLwO7aIPc1yBKlKdpqbwqpjs/1/TEk2GtjmLNDUGIH3R60SMcJXxDuh
yll/f+/cHUAj0kTMpQPegq57+pNVQta3XLPXUlyDcq8W1pbCZyW81978+C1oW44vwd/rIXlBsMiy
7GpuIhCItz0AyryonZAALZpIwHAk7zjH1WC/49V0JlClhtqlm+a+GJg87b0a9o2+6h1Vuzh8iIqS
LBVIWMeg5YMO5hpowDvWj50rxVadQbDA5YK3Cf+dtyO5I/doDpYM0MxriHmRlnAAvB/5NnTxyz0F
5nO92r8Hr1yKL6Gkiwt0ec04S8p0R4apP3ZJ51usYGqtxLnEU0SVRQrKq4B8D7/UPqyTeE7mL+9V
J8aP7z+V/7LsMsWzJFyd4o2CrT8Qry51IOtBmHvUQFVOHel6GSpO5tif7eRx9DeAW+caHxkkSVGY
vfc7Icbl4pRj7Baj8gUs3qGqaTrWR50xYxGJuRmKv1tMOJr8xfytxnnNAXNr7TXfHRqXyeEOUAbx
6jFWu2UmhZpNRGh1tbyBpFgi8rS1hEZN5HHzb7eMs0EhaGnyFZe9IXRB2swHeoMskUI5EZARSrzv
XaRvOHMaeyFGc21i1cyTtC8H3H61x4pS/Agk5Cwi4Vtvlfg1m0uI4Nm1z1bz08TbiB68r/1egUbT
KmplSHbnp1yAEM9lei9DBhT3THUKvX/slni/l6sDqCrWGjwYi1wxhups7q4bkXpzcwSAkZ5nIC3z
DZBkD/C2EfGAqGSe2MD6DKCHPUOWudMrl6BVllYT0qaRYlHWwt8qidoKQb6UybYC6k7IwJp+2WDj
Avo17OmbvxDL4RKWBEzAVkH+t47Jzk94Xv8Ezy6UYedNkkaRA5/pU17ThX45wY3leDPcMdw7veBr
T749Bjj+BGg4ut/SesWGoBvdgLVerjlY1kpEqMO0bgZv+acbKjD+tt0qfgqbAgAHTFflUXfjhVvm
Cw17cGUp/oOyGIc+TNArbfsuI/9/wH5azFZ2U97e5V14paN0EFLoLmxJYp1sO77bE5Oaf0LetJ8F
zbFADdakb+vWy5+Om1Yz3JlifhH7YxYXsuG4m7UkIrDOn3BIvNpp+lx4EknFurXsNC8ip+Ghd+8A
sU4P32AhuI3BFsXQfo8fr+vPyhD1+qCKCRxeHW4e10zBEwSHCLhL5u6AVND/VB+BhYSogG/8v64s
8HcU7Ij3T0k+MuPuNwwqodALsBbfRero0fiof7eEbx4eRwH+0FJ9yYNOwQ7sL+MC2TpeFKKZsXZ8
3zYFKgaaFi4qT8VeuHikyaPccJ3+oPzAPfWboXqH5nhXnSmMf3DRzgF+QYtoEBB7nD+/efOt8vdj
mPe5huz3C9fhgA4Hl8+DiHAkOOzikz1ES+oTg7moOUO8RfrEajdoBfD5do9mgAKjQ18KpqjAvqvp
NA0lBTPno5NkZLuBj4eeKl1cFLD3m151g9agemQs9xHYqt07YTm9Lb7x1JcKY3ooFwaGS4BFaehb
GOrH48JVS9WInAEjSI115oWuGfUYn40eZMxJ/xcLjsjoTT8/anjg0gtXfxjAEQaS+SKwaCFScz9u
r9t0EG1PDnYMnwV8nBso+4PkLmUPaxIcTmoEBEP2AZpyWh3Pf5j8iYosgaqQ7vTUpHMG4w2Bpiq1
OOAhi5/MioCxsSn/I7m3WpsMLxZcTIc3xqtwguclNYmIcSGjFwIYYndsdpk5NxS0lk/sb4g/H/2i
Z28wSVWuJqsVYyFOwwwaeImLT1AgsMobBvbfFiUnlW3M9dpep+Y2BmccuTYwWbADlQMVpvcwU8rI
HbaucThbbX+sgxsJmWkyxIQAK31RHXwbH/cqXcvE3TAtR5Hfthl7CnoMOTdFeIOKLF8Dxl3/3UJ/
ziMT/88skBVarGEC7wfmkIalMzBZwyHmslOC2dJP72JzzloHXPlrD0AS7cdCFf8QcZtxzAGaEyM2
HpLlT/uuc/6HoAFzxXqSD3wJPOMHLKErzxQnPqm9y9Qfkw/yqKvJS7vFB4Qy7QxdoSxxLV0b66ce
f/ex0RlOm2uGLtow61jnu0n9vhYZ8MeXh4Al3eJ/PzWPhV2USqp3RgNF9g3NAbEZUbtGVIdKaZoi
n8OXC5FqcaAsmYzWTjonCbdo6NUiRK2X74xDRuuSdcoQyj9cucaa5Gif0RSrpQtkivRxrUwvyZvU
BYJMO0KwRvcKSKbBP1/+Lwo4YqrsEMXs+02OCXiI9OQQFhWVXbZOPmfsZNRv6eEEXv5cNW+jHfhJ
mi5P/lKMuCggmEwOjSaSVGuxd+XHRIck0TwPUqGF7hEWM3L9NFkMTEpJu2hSXPNkwCAzjCgIVTjW
CJQr/v9eRQPJWJEQlhfwPmY+AOPFcSdbUtEnZSivHfHkBOJRMgHFVtf/7ht6kED3tJdZ6t9ifOsd
HOMf4NtGenxglRfGdCTl51nBAY1yAO1rdh3XIadmBBmkueIP2sJQ9nPDhVEm3p3T/+PTo6FDweDv
VWrVtpkt+tN8fcsvCsk3pOROrKAQKNgxZrhaSrWEMSz3SWYff5lQb0Y0cVC+D7EjxoRUOjNXi+QE
FjVfdI8RMy3/Pqxj8KlR1njvybvGr992IqiWPAncmWXFf0G2CsH8+onOVfCgt0De+m35O5CjyNQO
o8rBi6XtOX6XIh5z4h0jxwQgoIqB5hwum/N3LPHb36IIkuFj2Ai5gEFm/nN/k0xIzmqts1u02l+C
Io0g6CQx1JW4yBdvA+ZEZzM1t9Qc0UDA/LeSbrwATDt+ZrknaNDBmq/A+FRX/GsC0DQd3bSQAmen
vonaoQKbF+BnIs3CdzbtJ7pAU92vP8+ZZfPtnyfdRJmPb/021ITdZGs7RMls7USXKLxgDdO2jRUS
KCGNjdceYXLGbSJyMPGOeLf5tZlL0MBvrQwI50YTRUubO0Smpwv3DBD7b7yKPY9S3FSeu+mBmCSr
XFE5egPGDtSFlXD7rOiLyth/oB6BlorF7WWBWcAGQ+TrVcPfquflbvqpEpMR0zPRx0RZj1Q/0Rzv
50pI/46TRHzYEmlns9PQz9OsBF2TKCP33mV9kG45DjzFIvjMZaAaudOu35/Ink2g7Vs+jT2jv7zV
LyOrA7yafuatQoeVkwMTnxGBCd2TVX2zlcQC4gTCHj1+zOzbLwKdzANqePixTihoc9mIpDvVoHJl
jwiJ2GmMjo+TvvotOZqzo77Zi89BYj6D/fqMszS7BohRpjJyRc+eL2XYcByCW0miVxF/N2tNr9vg
IhiE5YG82yH0CFTEvbkHl9KcIyO3ckPDyDHV3n82+xev6Tg/fFu5MHLmAW4ju14Um5c/y4fXxcad
i42J9lW96wFZ8wHnfmFNCSocBR9ux/Lz26Rb9sd41ENFyMEbrawl0T7yJLHA5lLZPjOhmVLQBiz1
Lv2Wcn2yAtkF03WIzDUUTh8CPFiqaazt5uGhesFPCibR6m7E+NFLmv5/JzQLk1oKLI23B5HxpFWV
2HJJFAho8mm5im0IG9f7s3uebI3U4teV62EeYKL6xrln4JtbEToL/3ccjVhqRf6SXP7WAuz5bSCB
5KzxzO+jxQCcD/c8pHHRXSPL8tTNynlxTKNi39zgkREzjzlr0wI+Zn0q2c5pEGhLcAGpYeP8lwTo
UPbnYgBOYrrL+ooyaTDKThz+7H3whUWFrCDoUOBh7eqh22v32vD/Od1cwiQuRCt/KmA7kY5hm+Kj
ESRFayccRqXimBKDFInhqRugWS23zoFPevQsoMNQMIZKDbZ6VSa57SYsM2IgOv1RvIDNI0aQnDSm
GFv8UH7+UYZC0EhEgj2kmpDlNviy3cMBa8uTZr6qnNHNCyshqSAIDi8v/66rdkt1xNc842Nj+pic
JOEp/P4n222iW7GwBzd1SLRDos17W3yIahhbR1SMPXJLpgq+EqFPkMGrowOvNFGV3P+SU1vH12F5
PTlj58f54x7FS8kHGJEHuq4Iqgjf9LRpjYQD/Mcsu/FxzKvIHXon2tpyf8Sd/frGRL9/eFwPM3c0
iKNpNMU0zmSwpdayGRV5b1+pobUzd8xmoc+C9a+UlcjP2OqXa9sR4hnqF5JwMmMl9k/S6XCtPDcj
AraVx4QXBhLG6OAoc0SxM1s4Az9Mz7Q6pa41c6cEgyNi5HBfQOK+BU5Z09a/ZGJSJIco4g25n5+o
6D0DVpNzP8KNiiU7g/GcxLj2TI+a85IPwNj/eDilXDXqGw53mdGKBsH5PQrsYfjEZqMRmh6Ji1S2
+wVpagxcfZMTE8PSA5o5bNsxddx2bSSavylpAmzSXpzxvvlFglGtUyUuzzP+djoDe2i8IZ4FRVzj
l88A6rT/ruBH3PVbdqcoAaukrOIJ4ueBqC0VULiirFW5jcWTBn8FFJBCvz14NGGduNCP5PcxD70C
48DdfK6XMZ25ETS2Ef+e2bhLrNP6gYjUAxZpjImz0zsjQS/MguqaUFdFDOCr9CxWnouUWn94Y9jv
bHn8NZ8t799NOttd6WwmtJzZBUBk7mOklDU7HbBEntCX0k6boCFk2zVXVmx8dXqrRstnTX53Isea
sCOlZFyLeoFt8GJyQYMlmERZXaYV5cdhcLrXXCnKf5Hmrc7FjNLLOh67IDjqTQbbszEp3sS/cJ3s
JB9sZ6TzBsCcL4TYmo/qUIoLpw5M2mnU0WAog4c6VM3oBhAXIWbKIoHiuqE1HO9zpQg+dHZotusy
YgxtvSrK45E13bqPFZTDaz8uhQaf/4IdoOVGuLxvPlwVRnuuKenuPW3lLEVoS1ciurnlUinXy2cu
jzTimsvsIlOgwx2QDFdep04GEoElY7OFjPsup3gFT0J27DoFezPSNpMUGksOBX5ZkOPA5CLTsnJ3
L8n5swEx9mUYQu3sY2pe0IG3d2KCHGgLV6lCz+VpgwDKm3hfNRt3AlfAC7JOSoso3kBM2RUeKK2P
B5juDkiJpYrFYvPnbgsGMFOLsULzkWvveawzcn0erOXTwNrdMcSmRPawffwXcGS/e7Imjz5bdOBQ
DH2PF8XRaho6F9anUKChS69sTcc3TNMnicAo4cVkMMhhs5Etzn/c2m9PPi6a6gS8nnRcyfpIOFPH
DU42YFpYeikkRWh6jIxy30si43SDjCCYYq3eaZfuEql+acHFd2yhq4xfvsfKq/655wWdeGWXvqBj
OyJZhieTt9115CA9ah3TkX2StCZFPNsf+bA2LZ0AokIs+dyfAi13AH/KqT6WFJNQwe/IwZDfpA3N
9B1fcum201c/EywwPyqNm2xlxmwTFhT17CC+b7Csh0u6OjRF9KAzxGYXQYVYlUShKzoxSzyOB4Ry
lC5bbqoZ7AdeF7vepgLCwdLCpF7iqzfT0PCxjsN8U0BOPqqGeUsoQ48hMDvouxMEeeKxzqAIpQpv
Il6KKrWLguSKLG+vR/n4VX/MSf3yIkkHhokx8iymzTDoXBSbg7DW0g2pv6iTT/ejHiZ5yYg4Jny7
G+0q4fsySEOl8Lzc7WS+u66nPJFm3Feejx1xMM6YxU0uFzDZkMMiL07mYtXzQGpssC8nvGBJ3qS/
SL4egZ1IaEOP/2AnQG9yA5cZtpr6WrGl0Yam9n2GId4UyHEIHtVtYandTjcVzsWr/vKIKQCjLm1K
oHsLDYHEuatRUlOJ06Le9kYlxbCtBUmW7Q8BOt5Bm9L02W/kjzEUseJ1iRURZ/WVIccDU8mmHdGG
sbwndrgMN/d/xcqxNrgtLmQNSwwwjCSuVDu4BvQEaboMzManTO/KztcryR/BzrgUCt4tbdRjV2QD
XnAyKuT6XR7BRQ1AwiCxRdS1osrQK+GZ7lvbx0Rwcly6FWqqYnVB7zq0tdH4VtIlDvdUvlJ7YhFI
oyI1ZDj1C9czZ6gT57ou8Jp5+Gy9VMtDj5seSHKEAAV2DVOUGj5c8Ko0TN+OTYI9G9t6KCFD56Gu
J4YuZp2H/W3uklGY1H5lZCIS+bQWnTB5418Udzusj8NoFpPJyXnpxQln2XOIiFf25yQfcSvGVdxk
j+9zRKSeo7eg5jr7xv3Qr9nUCtUPGiuV+bd0pyOl1eG05IwjRM2lnehfkNPsRosw3diP15QnMF8t
VwcDjyqpL4pB6wTBnsmueCO9HAdpCklEl3MmvoFAeGejpyzWXRW28c3z5niapq7vXJ75KJ4f7+KW
+Bq+vF8r8fCr9wJ4qUV6R9pqC6IEjtqyTGa8l9teIu4g5zvi/n1IfA5npyS7lXtPT1WdMKF0NRIo
Epz0/BClq8tdlef2fVqnOSX1i4Fxd+OgkDfYnXyeOGG6Gs0iEtdMoKIQY4BjM5JX7lRKJNO2nKn3
riuTFBQOs7s1PxGkHTlR/1f1eN9XrT/ueij4hiX7rCP00ar7BlskuzgIteR8XgbQizHbT3nJVoPL
DJSC9wxoY8I9z6lB01hclni9TzPQkSaabPD62BUFToxK8swvQgBwL25Hq96yTdTSX4wl2hRRDHJu
5XzemZ2rnVA7y1K4jN5VU+AYvUxzJdOY7jzAaen/7oHPmL9hObclisIIfSGZcRydKaM8hMAZP6gI
ig0IDmGvsjaF/zUcwCTnI0623pKoYhLjlirmob7ZYlH6tikFVwfOs/P9vRmsXkLrtwpKKV9xhPvU
4QVpMNLFTf0mSPsViexnK4yxBRsdCaeVohbjyDSHt23M1wo/6zlywlCQkeRTp+EcE+C2UjIpd+SA
eaB8qZwpfdmc9DAshMjcw/LxmKORCGj4CuhAAgNmAy1prf0ExT0pyL+1s1l+xt87MpojWFSs2OQO
MlDyeDqBFpHXC3OQxyzoEHeVkfLskjWtdpQ/YkSui34FGnllWDbAXwuBdVsWzm4mltCfv29DlzKL
DkQegqfUQX+oA6/ylKtn9mnekJ19OyJDrSd3i9/ynGs03X6B35vKx40iZVvNKpdK4xchbLePvHP0
4dqAwdPbFA3LqsZ/6EIgfBlJZY6a/G94+JMnJWRBSLSsZPd6lJ35Kyd5P709cEDBJQlwEFJ9kbbk
1T0+S33WvIY+mCmBQLUhCSJLLpqVlxyyNtJb2ZNRO1/alCndHGAF55UseBHtwwy0HoNNFXSIWuKd
3+88oQwYI8j7zkEzQGGbA9IrXy2/ZxsW4FT0asDEpCDLhypOkY8sQkNleensWIp7poIF04EK7r8T
OcEsIaOss4RTDgXZ7s2y/WQ9UmiOPdCEwEzlhHHi2V65ZE+hwKQXMO2IOLHrUUBKXq0ahFpvAQjo
K2q5c94NXAhdxwqFJUUKQ+sB5VQ9JhUIM6HEVOS+HrrNN3FP1ymmE0IA2V4NTIynz45i61Tv+gRv
OYlJOLtnxW9sBf7Co0UpsLOA/wtt18F7xCyGGVoZL/5lU1jtPbfr9GJ90B4H3OZI1keu6KWF9HAn
6iPODSI0tnFON3j+EkS1LgC0rEk+dbTURre2W0cBHlWl2eHm9TWk184qwDczviKryy7B06dkNq0T
L/PfgcGZS4RtpAJp/l086XwcbVs1eD3gXjEW6FK2dXaC/I0nP9BBZ1wbvHlUs9oTrtTre7rNAnIu
AJgrJDwKULZWDb/Xt5aBnPQCkEBV+mHWTPWgYVrcLvujOhj8iN1Io1wUi662NFIvOyn3AKzBjbW3
mc5MCkf+IyHJvHd9sDT0C5eOhIm5m+PoyCysEmEMUneBUyutqaRaA7dTHEXpEjKQHguvilisaaUd
6Ir+TZZjGqqavEXVv8He1PgC831GMNXANHpHC3oRlhR1W2ybZ/00hi8YJo9OyZLeam26LwJLtruO
EBgd3qK7HdAxMqrAJuTj0fleTCrPKZ9U4ZubgOzJ5XMKSJttob1K5GUiiIe4NFnRShCCOUaYijsl
i10ey9I+A+zqQJXrtC7AVUti2wIR2Gm2KfOVtUTKGnNG/WwlYmaElf26819sclLmR4eYSqx9BmCj
uSCy5If9aXs1UzVtsDohwFX2TzL90f7/+crpdx8nELDUyl+cm2kpVMoOrSzPyeW46+M3GXgKoJnx
nF3ONSwJ5OMkgU8rY1fRuGSzR5LmMk2Sam4MeBP1teoIx97YbFNSpxh52oPQUIVoSM9ILHa4KYlp
tE5Mbm2rCAXq42Lpm1uFiEZn1VC+Rik8WllM9E6Yj2rmqpKSiYYvo1BjGUzWIBa375fqM+JjOdmp
vIlHok6EA0W58VcX/YLLe4kXAh0OfSFtnZ+NFiQpQn6WJmPeCbov7cXz7BYuWv4nt4p9qZ79Sr+Q
Ma/t5zUtPvktoTquv7mvthws9bf4N2HDczlOIQJ9mYOSSsNZNG7BYm1EjYsEG3eBtup8iWYKQS/q
6yL4WYKxaIY1o+NlmAkGUj+CZ/+xZtcJUal97Lq5JyK5Xyd4bOGKIXJzXc2erQI0gcOuXCWD9GHr
ptxS/dJIwQHSjk6JxMKgZtyO9OLZNpUZV3YTk9RWmaVvVVUbenzdRpmp3obmGGDjwwxy3xmpq5Bq
dYFXGNggmkWmz/4btsInNf4Xl80ubzgQKV6VF3FAkiDrc+lrXyGzMAScN2AhqHPMvrIta5BGjD2A
bDNkuqES74QqNLPEy+A0s/gH2OUYgaJWnPt7+Zl2MB+qIbDTXSfOzBGV0MUJvyAqTOJPqZinm4cS
1kDX0Ah9vaZl17SwuNPTDOrLEKJ8WTPxND66aWej7wjlIvB/uy/UXOmpsPnPZVuqhWSad81djj4E
UtdS2EJkaIFuDf19aJDUFnQrtOSkgf6awaqFE66F7AX+9ASbwR2EQldWkeREXKXgZyv7YWwiCJbD
7VhWeaH0MxeuURvo7KxEq+RwFvOGbqBHxAFjyXz3EQ2BYnvW3A8zTD2i4zhlFneSVMtrqMlaDoG+
XJCERWT4tzCy9fUx7PqYsd01E4FosEuToItXRS2BByVN583099ykHy3eWQmaGGWv0xeXGdYYlLYQ
6R/RlydULxFtDg84TIXi4PApMHckmo4yn9wXwsowFJYer1XFZ6PO9XSxQjIAnTrtYZFUY7VlbA6T
KvaGYr+NCoXhHBRaF9ViflegM2oEccf35rtduH15aBliCqks6upYvs0nQR8tYkaUfdFp0hp2PC/Q
RCE74vzL3DsT8NN3zTmUviq46EDZYDKIJQgoWPVV8oUgfXxakYRPGpRqV+iNNXDRaz5msMrYVG0T
rpI+qq7MfMCFyVzA0fMDweV7IHly5w9s3UUTHC8NHI4JJuI1oW0ngTQGpgrsu79gEi1V7F4J9s7X
cDcw7YMTsmTbLmywK6eU/vqEn7lA+Qu/BGUFEHOV0dncXYawLCxstRJQPpXYFjM5NlQ0dZ6Q8Xb5
YFgHPoTzfiBLJli39rPcSrQIikM/4efLkGNG2POz2xfUZFX8YM7qACaJVkuXFSqnKg/BPLgFuJv4
bt5jA+7Z4PB0I+Lgl5PKn6ZJ2bRjnzyofMXv3QNu2QaOpekF3C9DnqiKH8EoAqkSo4oA9a9pt+DY
mriA2ZfFJ8RSfo/zmLIg8PvvkQM07uPU31yTIlVpQdfKhVGE4kc1sNkaLZ+5LTsXsw9lBPIlSCxX
V/nFc374wsv/prumzY6pvyovqCGDLUDL//05jEKO0gBEdIsTiUXLbSv+uLe06+ltlf9DCIeXAQQj
jfQCMKUF5oNcZKDZSRFU7VA4buwrGTJQadOntA9/9arW0M6gprZA4IgDONAAMUogCzCfpbo6N2mk
Dab1ElfXt9AJAy6H3TcO0ncvICIytroHFVyQ7CXH2oQlY7De576zb/d52SiX3TSyRrSmS6LSDwGr
i6ja/cGAtT4kT4f0wezj16YvB+pm4PyYlkjY5k0Fnha/Tdd4c55Mpwtbz/wEB6UWd1xYGPAFLXPZ
Opj7IUrkBUvt2MlPrGpUicG9eqN/aCzY5h7fFN764FwnL+/yPPrbnM5qwkImsf2jJ/W0U54YXw+Y
GGzLNQYJXbOpTcXLwLaL9gyivVyiERWRQSA2TjLOwvWOu8ZuHoXoJphSS5qraxIA1XqkXqRIOS7g
ls/w/bJYViOq1DpNgNIDCQV+Gd5b/k6/XZjVBaTadQKSl1daGflTCxiaQhQfrT02eR42ZLDGIifX
u4t2W2lx5GhORuvwv5k7rms155fiJEtOFN5y9pONwsuwYzBLSWp4TgR/oaPcsl34lJFVZe4ZIvcB
WuFAQn9KdXmaDPDDeM+AiXO9MOrCjQvE9numYyUVLfaNN8p2qfBUDQz0MaqYFgi2fiBy9J1MbtQ6
5pkInyN6ru0JeZokkF4JQ6atRhfkfW3DV9ugkxQARJEr8ArMP/ZRHNb0mmeVzfQsP9tu2bo5XhfV
48Z8Kb9QZSm58V0tPybo4gu0bbO7vcjTFpY6pR13Mm+dJM7g6AQhVDlH+jjR2Vf9VqJErKQcvQ7n
ZWlcjL7D8/04izleP8hB5WylG3RB55lsMQcfSX8XeSQQiu76aM3GF3BhdJJTJBG0sm6yMSBxihZb
0efLuy4P/whwiFPRAOArTltPlwNgTPAQvTcRjQSIQRLlgRrXov5k8jnVXQW62DkJYOsaVxZekpQF
1stNVAFb5Ct+zyfIsqZR/G9OVuhR7kwwmTGtaMoH5COq0vnDi40d7ZZKWw0yrFIrFUr/gDblmef4
EcDpAPlrL7bHB0OGp3fkzw2RKmgfL/32OE3nGtnUD6GFUB7yy+B+oc1S1Dpsz4hdac+koc4NLSF7
me9epnjGGXwW52kHxuJHuxfK6HBxEZWkGlLjeddP7dVJ3nvG3cZzanNsdE2yBRlHWUJsI58J5tYL
CyecWR7bQT2ZbnfRAU4BykNUAMh4rJx6R83iDdguOcQVTtc3keS6jWU2cpK4QKA2OIqVfNvI+5gU
UCl7c7BRjbahHs/gJGVOnGquJC93fDiOEimOMUj1e5r22fafFahdkSCd0pnX5iFvjW9msiBxG5Iw
OOB9s2R8hnvoIMAm+Eu44RzNlAqnjh8B4DKXJ623J8wii4KeXMUklVHAXSTESWWf1ubYommJbOuC
0Hc9EVbYY32IeoKzXwNnbN7/zAPYknRNmoulf+lh63ELAi5wrPnv8J7eDwE1UKhXJ4n4bSWGJmCx
gO8cR/az4dXAm5UEiGtnojU2bk2heTgRbtfWFlRNDol9sKn/velrTf7EqIar1gYO/I0LQb8JvqFU
UIG5bxPieBzFz+C5dvMjAH8cvkZ/aQbYhyrGPX+S31WMQNN7g7Kqprm0KkiYyslXVUHtQppl7MYQ
WtLT/26dnZeQ7j/gUlx5QBSzbxQAlb0xzueiD5Lz/O1isa7Qn7BemkWg10wfxV4PALma/6OjpID+
/TRaOm8FOzfd1Yg85UAGrpbvZWzi1ePt83VrttkYI1VhnU1lWtsOpUaObajogp2MeTQu1WDvbgmj
3BPD6joRY+TjjFkGsSI3RlYsKCQzJ5AAXn+kgKLFIYRpN5oKQHt//ECeS8ujLJ/elgnwK2Ifwx/9
Qj5Ts07IWsECPiLbEZsmhjJTczmlgY28NmaW0387PzEEBpP0PZqNHj2p8alOoediGKCcG45pkZ2l
h2iTW9KaV28eLfN5lI2wlYbd3u7/ExpG0Mk4pX6+w/s903wS2qOkRW1a1mhn5oY/O5Q4WEdi+CTH
X2XlXxc0TPhCVg5B8mgsOjQdy+XB+5XXcsdV07M5a4ShsT421caVFQ//KSiiW93mWI7DNclUHEtg
xoUlWtpzHd/Rw4of3n8y0fS6/M47odaQr8P20v5uQslvhFR8ckDFtwJGQe/BxGM1hwOCC24oX7uB
FSHxrTW7KP+sUvL84iyz3MHdOYnV/q/R4pd6EXuBMcZpHxhCcJRk8ILq/qKGPsVqeuhiU0f6p4LD
D3dJLDxL00kl6BKPMOwQtbIlkMLpx1U42uVG5vwmXrBHNKpAykwDzgamYkwzgrW0VNEM4LhS0JOs
ojC9cSYO0e84A4MOJlkge0ylNWFNR0PJOo3XI00AcZGzRvvW1vkU/7c3Eye6FVA2Km1pseEKxIs9
thKTyciXa8ftFg+qglw0a+Tb4yGtQ49wgJsozM7PteaC6MDQJgRWE4zShmBY5fK/4ian6JPW8MKe
40oVsrjiWmW7TELUgyLnQeqBBS7gCOQkorfEIn+0P5BEHQ3CgnX8Lhz79zDtD1IzRfRrZ0GR+Nf6
M0d6Vmi+fcnmQSob84CMgEb9A54xgUI4hKUl0JpC2co0OGyFBm5sMeYEgqomNrDTiJcD8iypMfSS
lm42dRCkX9ILraLOe3PYda9DFo1z5aA8Kc7aGxl3SKpgRkOrvg/ph9vTlcVuBOi8as+/KEkcD4/K
12wbRDLCjXBaSHDD7qL14pRjRu1Kr3vnuXXoapyylkP4KIj3m35EnTKGrGjJ30zjhoiKZInvo/3v
x0KeLQk1UrPws6iDrDxqvLSEWY/POyEleCMaXP8QoVdLRYM9SDV+O2q+B6dj2fp2xi/kV1GbmcG6
FmGeChyP25HToBI8k3UAludhwOyKutMzgGXvmeaJLS+tXIfDQNBnnfP6TRxuFeH/ueYQL17sB2mS
OX0jR1v/3Jtm65X966TpGYLOJ92kUPr+l2os3IYHdN0MHDU4MryCgjwQIugzME2YrqRM5gFlJ4L5
9Rt0NKYe4/c3yKRG5CQ9uKwhXl3UzU5LHSYC5vLqLJ5aVH23M4jnFyitPWJDKS4om/lNcpPuKdyl
NO69K8Mqd02tMF7eSW+WQ0orMLh82SCG74iolxca/UfWwC+jIZIWH3Kv+k0XG1kf196Q5HbYtnD5
YHQV5chi9khVoMnjTs5d0BD00iLTTsSUfyx2Tj5X7AykZHrMfNX5LvvoZeAqPOxe53IwLeLLtc3m
m9iTus7Z1yli7P/GU6Zza88hRz8T1uxZsVWjUF+zgKmuf51GzUmfsse9zZTNz/9A0g+xQ77Lpo3k
i8HSOPrtaBgaV38mjtdwnMWelnYWDMYkla8zCQl3crpMspWWB/NuDTl+0ZDV9qXgKOI8cVDHmegh
9NellEiV0ezgojmbTPXhvD1gkPhxbfhpaCnhalJnjEY3SOnYRKjp6JQSjL1wz5nG+mszhGfu1W7o
O3qz/ugJMqKiwezaOIeUu5FUFI47NDcgqRL5BHs9ig1Ns6U3Xib8f4wsPFbwrevoahkiDwdyhJWS
8kEJmp6iXWP3KZ14z+CSiQDPTSPOR0M8/9VxR1PWYlWH34HcdrFUp6OwWojzXbGjybJV2yOgiu3/
lKzHmVZrzUU8M9sCNm7dApIXnSO6b/hvtAtmU8YG4bbx2Kw+ZHPi2uYes1PHhx+xzZwSp5BrKBBo
ssQ50uWRKbz98fSyeQr0fXhf8MuvX+y1uYIZzcuS4j0cjfmK4kuAQdngapSBtoQxYaODKNgOusaa
ONxGgJBGb5o1edAtGeVyOqU0dhrx2rxzNkO/gcnzkJvV8DBkn2Sf7Wa9QlQJjPSAA4ezDBK6Bp9A
qfJ7HhnhCD71Wd+hX4L8VSyPTSkXYpAcS/W0RWujBbEo1tYrkW6eAI6jTyPIrspahV3CfZTRWEFQ
WEcVv+5qEmFSjSXgBYwKZEx5C8MH7MLZdJ2CrFkU9udEZyMSbEewhxijiVkXKEX1FRzrIriBh+Rg
M9VDdf3xVeRuEwlericj+ji6l2bQw7i/cBRInnyA7rtTY2vVY5lljnFW0gpzsYaJlHpaVxGmToYt
ta2bV4MU6jxNvGAGWzFTML6dDEo3XeqsgwTGhTb6FmasHkoPcSdBCwvCVh2GD06KEAzYE3p2G5Dj
/+NpkG/hQhYJVT1LRs5pxPLumZt3tjI2H0bR0rxq0yTrnErw3UwIgAhaov+117xsHRxfQYWIuLke
uA0lanPR3A7sPeGr3t3OcBpgCI1vH8Eu7htmgdSO0Jg8/Jk0a4PYKQ5pp4b8eiSipYAMa6DtTpuY
EhOm2VuCh3jbMLXLU6pkQgkqCFpuhisUcWscMikYLFL0zX97opiPxi4QvSF9vK1uwwOD6Qcmk/YD
kbOBeQMw0SI2coBYZ9xO8G1u9x7XrkjsurSGh8eGGIxHvVwMB6VjhRh1ixxirfMUy2fm7Z/6QzJg
pgj5yQOqdPFX8uwM0MyV58kdXxd9pEwbGSpk4lrxhx0BLy5zCFtlTmsIsRMcncQYULpdmfQsRyMD
kBdHjD3nysb9YrbViEcuaRifMxptbVV9Go+D3ccnrN97ilN0mZV00yaEiwIhDXFyUPGLcs6LTpnK
GwSa67g1k6LHPHFBAtiw5p/x4jlhh0nd6MmKJDoI2D0gkL0/fiWSH3+NbCjJIKPC0KxRdw53SPXj
xy+VW636dm4K1rGKb3WJWuf1uNH6MM0T8Ci8SCrSHQ3CoBPCM7jQGP4+oeCjd43ZtZgykoQ4GMq1
Gjn+qRyBofIN/2rMCPmpumkMsjKhl+kwLy9WywrvN7/F0jaPyRwowyzDfUuTLS7kSMR/oI5vw5us
gledg2cdpJ7/JRqkerN+Ru0NKtQnaKvKdoB4zBS2K5g1KB+0L0nqh3FVG4/NaZ1sLpb4ak9eDPrk
QHBEAYnSmljAbXp2K1uB0polwiful1b0AtAzqOFGKwp+bM/hpUVL0LZkJ6GImc04/nGNIYy7LBB8
FDMtw2aKIQDjTysD+aVysaCGw2zgRzh582shphM3/empUzQtH1/Ud9njgmgIAjg888lAbQh24WPI
z4umSC00DPIpMiGxzKyaolSClQj6gCL4D1qsR2e9iNNHiGEeO6Tf3YHHRrVHmv0BvyLQhYQb7qrW
XhUIV+C6J5fQYUwG/jav8qvXBfYgyEJSkvfxw5UkEfbsLS7NdEI3Qr0pkLIlQjoRggrfg6Jphm6b
HiAMiTprO3T13TAmi963EO2i7j3XILpnKMsRwc0uUZ0BCuoT1OiZ60LN7SSvTpdwyBTdTGSvyzJp
WI6n0J2yVgHm5HvzqJn4DL9TLWi4sIhOOVzPpHQZbcaRfG0gGHMeh67dR7Et7LrGBpv0DeOBDlXC
a7ODOovEgGqJ5ZjYNRNjzCoD54aG4Th4Ysh3GkjQRT6OQS6QZCBhrPeJIErJuYNIsEa/5WGh/+vo
8+KEhjeEobmuWn8q+mvkTvlf5uijNzcHjBPto42/K6o0aRl42ul0vvkoMTlB+hus1uyOSkkszfWj
JKPiQlkZYVesA5FCuAfPXFAc+k2e3KsRkL8gTkQgivQEP1NXG5cAQgz4DAqZ1wf2YanTmsk9NdTv
Yaymbh3RmsMavu56QaoUinIUlgy0aJHImZ/0ZHqo0dzf0SvNGOkLh6OwAd0Agkkl395MzfNBSRT3
A15cQpZ1Lp13IlZhQVlG0eEGmc3DnCgnpAqilspmKqVFMIC/unB1nXBelGEkfP3c/RBQv9rPQh9Z
FyjYHfk3xxc0autZpo7nV6mTpljvnmhSX9X/xo1BWhqpGn8HTHqo6YjRe8QG5s2kMRjdU7Pf6gwI
3pzYJhpdbHywgt0yAFnoAOM/HQTB/U6uxX3QGPUA4qeWdNXjTQQs9OgD22LV3MEBjLhlZqhudeFq
7FMBOPpMn/XaP75bH0D1L2iiZinfmudtlgdfQsQ5fDo/GgnjogwZkT2eYlIVV+9270YumnjcprZd
89zUbL4W00u5/MMCIdH5p26s3ouccZkHTbj0Co0+0QHdpb2S23P4g3CQSH1H77iSfgJWrVxTtsE7
lkIN6EmNMQSdPHyPKHqgaLj1f6akHtIME6ibyERMAUwi5fZWB07aWV5UrXEQKPFdA1wwbkC6Powh
WvCR77zR6fLydRHS/726zPw76ueeOaWupc1FWDhNIu3ogzsMZE1kro6I491R1WT1Y3br4joUBjtU
dIaLeyunr0LMmZeUy7gfbMBNiQTWPl0gCdMGTvIOvCGQvAlFtdzK2eMJ2kdznYkX2i+7t2TpSpXV
VDdTwqtt7KjqUmczRwBdPwMIa0AU19B8Y3VMeAWtB6yZyMSrXal6RpfplUKVEnH684rA2nw0ydmi
1pImdCl65LQaaaKOjmhaVN02cCz5etqsg6sOGNQ9EmphW5Ns+qxSY7Y7c6uSkyB+X+PrAojWmXL9
YHvwSJr+YMWADtHEM2+UYCEn/mbZcOCfJCaNxhvUVqgVGxrdYmY6z09uS2Nb/iCX4+0USSU6msG1
vehTt/dN68rQjd4mbqGfoWjyujDYL+xmAdWLCCufzAUbwlKER/FA6GmKpm6eyZv+Lccpvyu8U/RE
TKonoZ2F/B7jG9mgGUoavGDL6Cz1tD7XTmjeofc9/uWjAz4iqGC4uXqZZimwnRqHEYzEvqaCfTCK
qTVY1qboB9wOIZuYl5TXb29yTOWMnGNYESk0T+HpI/viy4yVlCLTrWkTSrGruzU4oauRBy4nauXM
K9Ojca0CIx40k/VK/n/BeEOsXiShVIh3lBGKMH9yj5B76RP6uDmPBaSsnkVV6+j/XlngBKOpt+WE
aFPVcl62gIZrWekbiwfeyum2940va/TINcp0sZStTCcAgfI+rLMy9GyiicqLsNcTSC8GW/0KlVOM
goH7tXh+NiYaPphEbPvZxzOQ2FX6XSHwWmIoq5xLe56Ed6/3g35cc00TaTHAa0xDz6NWJjFLBXmK
bQa+9tnIHDFJWhiVlUmyrQ3+1FvAWG/yXg0BfvCBqJfl9O1B47ijAbfMefFu0FCuW2SKRxqAdq8i
gZK8CshwLASkhnN9aT2kWfhM/Cf7ONZqAYZChGmSpWz7jBWEHDYV47NiFk28gqpsE/A2ccQLeKpJ
A04aA+ZMEchpa6LBrUzsJegkV4SSnJy+8Zqcr2bebOmgO3cbcbqIOD5dc/e+c1+nRONSAf3wYwJs
HkoIObJNJ3ZMd1jlvohpi7SqXV92PJ9COvZuHdyViCuA7mKVCy2eM/EN2hadul57UxM35V2sjgO+
LCUOVew/hRiwm7NzH3IapNgoTHUiTfMEg9byAYPWyDBkfB7kAapc3cQfy1R5/ReBgdlnCCF0FKnp
NokFLihGTfFENLcZaGe4EIoA55/C7m4WVwgWaXHyu0CfrefxywYlLC4/J77liLt8t0bjib0e6az5
6ElT7Cjs3wISJHMtrQi2eEW4905qdvg8W8k854y+O+Hi71k2Xj/hG9BD2V587rlsyexTxTmn9oN9
NfX7lfloWpKvo9mAIM6ynm+UFF6pjrXL/Q6fUTLlF8R8Psh0yI6oZQpbAR3POSfXa1Sk6zBFlZKd
I8C3ZG6TkTXiNIwyuoH/+xnGJO9UegSv01/J63cWvh+ZA+BAQ9gWc1CGoNIjyXcqRJg4T4hu9Qh9
K4vnmMDlv36poig8ap8hCtRv/FvI5ySgYH09EUdTWbmm//0GnJAuPnqm7BGtVivRpcM9z9mI0KPk
H8qz6+l40blKnl6Ua9IKxnCDEG2GxAuY5lqHJL10kFxPrR4kniN4ZgPvi0kgiK+/20dz8rH9h0LW
tsFPR0SZ0jvOOtKwNjBoqCOdhA7VK+9KPNDpIzPhB8gz+Rs14kkheV5/I3XabUJmFRgc0i8J/HMP
N+CG/iW7cfJuYvVYJUxdkVsD7ErSR9bRasEodQRwZjlFdoOpRCkECtpa5YVOmc5heC7KIrvFC9MW
27RfoZCtSgT90BjeO85tjgegLUQvzjFglzSSnzOv13iFLvbL1VrX495NqBV4lkBaqCewOVzPCWof
KAzNNZ4bYYYVecYY6mY+MHckwxbZMtkG6B+b2UfsF0O8rHzz5q59bOmBvuyjpctqdf919o2cji/3
d1uwowU9iJH+fdL7uf3MvYwOLoSLJl3mN5vGXqatRxgaP1qyvzGbQg3nhzjQRZwb5QfS9S1t/1N9
NG10Ik2YfZR9lkiMg8Bo9ou6JSH60hEkCvEaUQp+AbaLGg5M8er79HtfQZyRrd/dLCp3B7yhfoa/
Z1EN5wXrI/6GTmo2PH/yCyGn9iLY3W2FOYdCJpgyX068r59xLymNLzgtm2SoaJRgHEIXtNrG9Ad7
IQBZXVbysizc5AgagLMUq3YkX7eysGMDeF/3Yk6POYLDSBdVceX5arHfVciaHFASQ7HxPBx99TWO
S7vpctsSDLO+n0tS6QAocviG0gFwDCmTAS4QGGSk3/sMmC9HRsAyZxsePubwroUyMNowsJWWiUI5
2yjxNI3p7G/PQUng2yOw5GTIk44K1Xi0kbqtEFUPHyuFhhFAMT/UQcerzaDMTBPrC7DE4S+qpcXT
F6CdtlMzHdJsygoS9G8ascsSzisNGiZykV9F+YBK2Ro/O+1Nw1FvezL4lUG394ESSxjC1iColKm8
4yt22FcJ+nrVdWjbUOuBi0AGwMomlidvG2LWXxFZgbUjaRSy0p33fFhydRWaD0TxHQvG0mAhNwlF
SzSnyLo+wo9seeby9i2j07zyGdOoY6A142dYEjlHMFqqAYCzCYObbehveK9A5wIjZdMJThjOBH72
0C86M/S5mYaPnjmMThg9WDZXM2O5nx5lsjCpr5OVtFqzaLJvtxl5/puZj8nh2phY08BVPuNq/5CU
fyjOOuJYv7ZgbfPRU1IXQ3EV+GNRymsgIADT8k0M9LT+dbDSGHfH+70gM4rHLwS5lV2j7weXkCq3
M4wdf5qpfxVUFFzQV5Cf2oapnqVyBw/ASoVRdktWVOnxupvGuMJQ8usJYC2YDT7pM2DlZdWEB5ma
E/63yscPftStpRsTM9h1BX95YKNfoqfc5I38Rh054Pgd+kbNQ9ndsGrEnAVyeq8Je3z0RIqiRT90
NLQIfW+fFiuogDe4d7zlqWNJ8oF5q/DuTYJ62QwlDk+c7g1agO/PQCy8Ln515gV04WvUX47WLfMW
WIg9mSNWmBOVjem/hE7js/OV2riEQAB80h2VkovJ0bDJgtVJmrAHddKmnk0cDa0UUCHFsvctll2g
aIB0y+ehzqdeduH6ov42xatihcILXqturpMMBx/SPisaaYrOVaDwFM5RFpetXRrP+r2lufU3/1en
1BLYSphoVo8t/OYAF3vvvdCf+gvVSXPX/cMOctaPC/EwcuDL9lU58yh1D+TFstLdHJlMnnwV3qxZ
6ATpyo5ubbv9RxaUk1qGH6gecX7ncEG9gTCkn3EbSAdLT73Hwtvm1P/8PIQnI/dTFERNv6RIQnpe
RgE9PWSItJuqzok16uq2klm3qgLsTeH78BV6KzxNkWiZtnj6Dzlw2jObNYL+39yl5LYcPUchcepD
fqGTDmv0FHAE2jRRxiBlk58JtNOnmz4Z7mNrfqfxsWShmIYNOvmfOC+tHwD+AklfDLwIj3wJQdYj
lHT4KzvpustMEXOzwbRGZtNvKY7xrShjNvGBymt+4Ws0BwwXanBZ1Vv45XopINUYrr+JD+L0nAeq
yqZQILE7cbJ7rFinynaU8AUHdRfapwEGBtLhYPv2959h18usNw2xIuSEmnRPl2wOloVdeAOkI8+W
Ojo5im1xVaZ3hV728FmhsGpwNpLQXx53F9YM96lwbCbjYtMDxehrSn0d083O7e0BFLt4DycWIop+
3UwH4orH8AXGbUKJ9LyTPg0AMUWIN8BynUyajms/sCqIgvngvQMZ2Cd4wf7s9D4bS9Tth0Y+EtmE
m+mFoB7CbpacEC0CjM4TL6iHiD2vvJLR/xWcqrvhpnABsHEaS6suzPshCSpCMHewN4nKOYBRPbun
cbzMws88g8aL3QVSPIp6XCElCYuu/6N/mJj7Z6a8KbHA93KS10kjFGKu/CrXGmEaIEcvd7oOVvP5
nLTmWGdUfcXWXWtzl3pzQG2KIkJCW+W9B03xspeNCd6qfe3f8cfo2mYBWpAJ2oKnAUCP5tprdGY6
2zBe3WT4HoGLSd9SgJHsNujiePAxhUpTV4oUNQ2crPSU4yHtWpQTKZ7iQM9POEPOfHLLGuAFRRpO
kAX4EVAKu37Y6NRN+p2nuJqttTyJq5b1U390D2XW8UqXW7Cg6bV7UlqnYb/gmHCAmv+nUOwSk0+d
+xrUm3DBw98atky5Z3mvNNoF6TOf2tkt7PriPiU0I5mfOaLdpuLLuHszZ3VZaNm9wZ6OWxZXBUDy
lnVIqNe0c/jXI/xxCvZdG/8MEhkHxUS0lhZQLUFxyfRYTrnjpkrT/i4YREQoPUdR0CunOv2UjkuF
626iLmtnk06rz2DL00h8GOWGrNin9fEo/x7FTi5m2GU7tCQzspPTPTOYeFh60AkPwujaEMP+0vAr
kOVwyxwb+j3b5vYjnGnrxQUTGLehl3RjzUwp2hfhaATmtfnB5W1OEsuQmJmxe7b53GwC393GING8
XGg85zF7uvoQQSx+qZYrqQYyVlzltlWZioDQdkl0f8UFmWXoYO+mAspCXpzwalTdOwk/xan8xkrU
8fECCksyOOl9q/ZeyJIwe4+SNosnKRRwrVd8M9qyR1gEJ2QQqIwO1qEjINO16tqUmGaxZO7Nk2GR
3+nCxo49QWKKt83fBS8FAog4Zp3rvv72Ci4aBwo0lDXu2NjUFp4ZSwlXSazvA26kOSdTlD0YPrOQ
9/8k5X42g2JKrmdnTQ8ETAit13k6OCn8/PFfxoGryKs1c3X8UbVqKV3lw+b4FeU1+pO9QEj2MPc2
Z0YNGxRPkyMjANFiiAeoCPXOLYEf+VulKxRTjTI1jJT+DGJXoGOdiz1QTA90YRBeXDqVrPMmsvcY
WGNUYCdFyKQBK715M3M1nK0TJpK7FVJESG0CBM5pheBKw7b67v+nk7l9Mt/NoKBfvBxlJNbtL32+
XOOhUWtUdXo2+aYNGAtHiWbGmMgLWvhdVWkUP5rsWAhirkPwAAWPTy0wIReloe2XssVQpARdyFK5
ynw16+jWqgMb/qYfXszMaP0l6Ufi3q6/C94wcYn4xtrW8Xuk9n12b6MxFb+3YdqVpmTQO9xjidsg
kgy7+QRSN0vIRKiXBngY+bd2TfJPrOTwVAOR7OeTI/Jmt6XKRX6IcnoIJEr5xiPA8yzQuFnh0D1X
ijnrORl9H9TxeeWMCbTCYsqewbHRBX5xvaPIYCJMIfyBxbkbm3VJAUSh/Ny3mPK/F6S39VvLMZzg
255Ahhwhjxai/m7T1pLgFEldw+Ki0eMVXhjTxMfiLOGGX1g2m9phTQ2ypxJ5Z0oS4Qxh1DFXO8Yn
CJbtiOJrtPWFg4m+sWUG+oiK6HoBfRktKDlIwa/OuiCXJAJbF4uSci3+oAUF05x8Z65cMreYGKdV
9icTTc1dSfnyIGs363XeSrEoyI4HGta0uzFBVvWn5vwtjvq+UnVILze8LK8xNAEU+yFkRulUZeT0
BMMsRzRJ5mo1sC+a/toZiGmXVZwQ90S/D64lk/Jz1I2Q4SfZkNK3+wybPJxqJBHVJ7rHShNWPkLp
ABeup+yc0tAFS6OTvuL+YnSPDMsvGwAlXz0mdMeMrU2uOfLrpEfH+qfSPQ1GJEv2Kfw1jIwBY0qs
WXTMIpFrWq8ayObV8BruZm/qoKDmUikYqsl9sQSA8OZe5kSehfc1+JOQRlx5Cx5axNCQ9qGucQts
XCAer/BINfx/FHJd7t73qYR6EskrWPNIeDKhp3cx/+Qc7ew+eo/hmTgXDmcb5JuMkJ8666gcbRrp
xHK3juS85kZNHuJlO77oJRjr+x1lY8DYYWIMDMtR4APIGbYSMhPcVaQcrQjXvtzg9GeajGRZvo9q
uLsZWjhERikqlGpRPhg4XfhwNYSnFd3g27CwIevUF2ASpYodLHldL7Io2u0XmbOkh3rD8QTVucl6
2X12mksRykI9Tfr6OZfNEF471HpgEO41MheHIugwjDSxi0H9u6UJDo/XD5mxgM0G3FskZ1+BmCc+
Smo2BYK/ikxp1FMzw9iCx42iRQW5xw7VzBS5QlCRU5XdKk9PMKK42A+519xvqYiKaX7rliOuUcQ2
9iAy9Ku6Ju5s0DKJvjw3mOLl/HubVkFGWuLpmwoLAO2eyQMMr5336McnbNo/6QU5TK8q4tdnAOsu
mL0bsKvkSUIGUJdZkfiiUnUlG/dhqrZNR3dGIRrvYPqgyL4MDfzee5Fh0eVGuk2BOjDHTOR3kR1n
VuVnn7JKvmIXYe3lsdREAzh4CAepd/Uc87IEUvJOxdzmt+aV8BizwHBF4EtfpjfU1VqBbTbM6GlN
+plEAXzllziZL1ou+V0S27i5jhR6qW6KAZaDEw6vjv1EFd+QtkxcZB50rTjm/3R5e+bIUJesI5Qq
FOtSe1BB1i91PcATmagBxNBIUGrBZdesEF2CcypuXms4ALmZiqoP5lp5u20h4EaDnzwRgtWNSJDa
emBM+VCggtVyokWJcdQXBj6P1GOlGUMeMVKq87qsxuRa7crx36DbLHvoejiiHU/N6cBTrWQF5P3B
VnOMbH81DXPVD755OoU4IEbOluEBP54yQQ+HhPqoMYSt7iTD2lasAc4pqX8D77PzEqYTEAm0pR06
rx4r2O7cw/kkzsGiHROVyDCXxgboXdVStJK0kZ3VUSEPGy2Eg3S18T7doOYNX4j1hajRejOMK+nT
RLi7hGJTGeUN08X0IyEJFylQldHpH04Hkp6K19Pa9z4MMTiUUuFAb5wP+aljsWSyAHh1VB9btdWz
wsfRfkCVNhe1+4KJ7KHr9Om55t4M1txxFpJ7E+6wx8vTOriwdtbcFmxTjTF2/ElO3ObXGngMoQC7
+M0WhMMWhWvIHuUnNgjiJpF+gL35rSIlv8pCOfORflNns6iVqTsoBp0j9D/exCmlxMOVzPHydUmT
MSAGmbPuIP4djle/tHqyHzQOKCnK/wneU8DNhBJ5rrlxrmJT6f20pOw1i8LLRx/D1kFkOBuGBPVq
nuciXUTULnXfCKWD1cHWTG33y24WnQUYWol/FATEd5ZKv4aLBN4vnGdPt4KvRnu6G10hDQtnkMLZ
SfDspJmSVet8F8iYCC74es4LN0zRrOjxS57G9Tn9ZTXxC523SxYd+bnRoQLs9rzvBgd8TO4g5Yo7
t+/3/fkQJaPG1GsC6PsnmKBC3QN7q5CIsrTFD8ktEQ5HiCu34p4hVIIYf5LPap6rWiMkPrEmf2rF
aB+SluSzfpED482EoV4E2LYSPE9DjJuI/vZYSilEzcWCLAbzBu+XJVbGCY8TyJOG3/QDXnKq75Oi
MW/BXIb/zUEb+iqbW6ieW2uftdENNgAprCVt7k45nS6K88ZmHsx8b5Mvw0Zqeu8ULVN56wyA1EzD
NRJ/Cj2VlNV3b9s4lY4Eqy8LPERhIXkdn/OSuJ1VY1wRhwAG4FpMRGQ0ifrRGoxlqEr9gc3E/VFT
XEklWUGjs8SoYm42XyJpeF9+3UbmpmaMZs8WfyToMYhw/qcJwS9YMxHeLpJub5InPJ8uPzJ34I2c
hBgxsRfOaelzPOQDoF/Jdkl6GYFsxviKxa7Wpm92H5VhyuVQgmYDOwJqsUzhRqMtcOkc7HWsaULN
IufKpIjcazO2oj3SwbCtndzmwH/zn//WdZ4blLNIiQqdPxofQretX361pkxE2+/ZYQSuGTfU7W1h
1euldZ/SxgwYYxpqw1i0zYN2Mc3eOIVgw8gdgQMc5TsFD5NKcb43pGZQcnP8dn02U6tdJaTUe6p3
a9d2W5jFdilNRlcg+Y4P3MCpRBTIaRtLu87/20RqVvW/n/AsDHVlEFhqXr2DB6hp4b6OL7Q4MuiS
hgL4k56l9tYvl1ICEsXnHd8nCz9dtrHVPJ8ogcUARXLyLn4h9TzgQ9LdXiS6uafM7B0tAGNiBajO
gDyqs6z9wlxnODTwO2dTaePegIw2ME94kWNb7241yizjyMMcLj+YrLPi0YiRcDq6oM3JyYGTo1pC
KVBHa0OoW8DLFc+NXxvBGwzsSmbaUjQNCtAOI9X9zpAqM4TCguxL441SG4wEcWYSgqk6NpyuHA8T
xTsY9rADOLfEWvIoHRYOiKz8aYG0KVwPmbgy5KA+HkE/3L0R3Z7w+09ljUOgbzmDWMLeLMR/9Lv7
XizpAmPUiVVNwCfRFO09xrh+DO0MhSprK24mBlUmNnAeeesDJHypV2v10qikeP1jMS2dEY5BK8OA
LTb8pUlCC6KZSw7WLo1iv+eoiz6ytTI5OISt9Od1RGX5buJOc4a1ssyqEIKdqeqDAATBHTHLDyRD
yh6blO2798Lgwzb0siKe1/lDS5ixpxbjvEFeC/KCfmqyP3e9bADEhwLaT3VAJR6IfsDkks0gn8Ta
iwH4tKtjkTl3/0CKiz6J6Q2/0WG/tpVquPJ1tJeY+Bozs77kj/v1+4AJmH3bFWP038+zb8N/OCJ1
fVjE/yb2Z5GhdkZfQ7W8/UgMcflQIT6vKRJDqnHztL+DySpILTYX2UJwR0O2lZGl7HAw8OBIvW4I
sqPjMzQz95sSdLbjZAUmQ4S3oD9uDnDnnXO+y1IsYyBbNqzvKlBsGgpsBbURE0DMlSk1BvP6hu1M
4/3Kfvtdyz3f2Sfht0VPS2Y1+42Xhf+HxLATqjbrTDcIfnRfTEUPToZjCvGnRv9IhqeZ04Rf7Jys
jwe8I8yr2R/OSi0iWbs87K3ElYtqt95a2R/jXDD+1/hgApMeXNFg9QtLwEMUCdFeL+lgpZPyrR3M
f6fIj4nXehW2GGQ//2XZDErPKobhQMvY3mZcnWhmZlf7JfgJxCLFTJ3VCJVonR1p2+ApPA4O7U7E
SMEG9tsOS2O2gQ0+3/W9ZH/MedbMaPHw96BneO74Oazaf3BdxuhilOTQljK2GBZo4d3gQ6baLERv
6JfThV/LSCanVsVy9OMnwrD37l0ZHYKiy2G0UsQ3nuCqfL1h8lMF4q5XQNUE+SngnknF2x5GDRld
NuP0ZhR5ymU0Boe1aM4dvu3u3X82gMqI85vNJZTeyuEeEUQWVMHR97naiAklljep+cro+DE8M8Bu
sC2hpR57ePWCiaSRSAU9zgyhbl58AHEwW1KWF58v4BJsFq7dkFCdm6ton4Z8n2WAEzuEi0BMwB+Y
+jJxtHGW/+fpLR/6MYdYdkAzl8U3Ii9zyPi3fRP+9z+8Dg/MRFHovwZTDa9HPrEAVVW7TvgGbxzz
jaMkG2qYFXU9/0x+5BLBD+DyQPp5BQFOYC/PvxANRpSiQ1VVdCXu00HuYMkMtg7QzTshWpfhTreq
6jebA7L1WVbfrac3e13sf4MA+PSZNVDtfCOXHdHgfd0d9ehq4APbrxuC0Hk41wm7lL/hXNjim/sk
Io3InZcK0JCVdcyMAt6f6cP0wj09lh4wRR2ZTLbi8Z+OvP7IEDLVRR3xtTu8RY5kCVTMZmRAw0pi
Hu+lcdQJHndmJ3Sj3O5cl5/WpifgIB0xv/fswG0+CjKregtME+6TY2FITp7/oMlX3vbyiRldp6lw
uMkALR1QLm6j3pqOiVWYIve9C6U5tuigTe7eJltEUSfOngMY1xdZQxsWMMNDECaKh0lGIMh2Wyev
dJOSWOq2xRkCiAguAqu2lkEoIHvpEUC7WO/+NCF857vvP89moq3wVCnyrkBmzNZAhfOof4q78SK4
JvvWJFd9Qbf+ZnKY5b0gQTOaTvbLjct40/vlzNilcZeAwW5Lbk5vMYyVmPLmLpQ0faHpO5ckqdRK
k0yk2rNZ4fncttNg29eopGD+gAVJD5dVl9maBosO0PIVnoGJBQLirZzeOqPFGJ5VOjhM5oB6lyDX
6jFyJNlRGikLWx/zHHowKpCPCg8IFJcF71e6DOOEUhTrY273AfE//j38URaNq9aB3puO3QiSmjCt
N+lVdfwSspGFjFFN7bK6l7qLarrR8cGr+trSg7nEq4RY6myWfPGTf1FAy1QrUNjpZFcmWon1UbdX
/OGTGMoiE76KiaThCtOISPTFyDnmz9MUCU/v/6FtgB60yQS6Y1AJHqashElmzGHNcdgdNdhaFxGQ
ubATxmYhznzieCpURqM7eYcxKSfzgDxE275uL63H9x8VCWQ+Rj3a1hRcxnYMxV9qLVqaCyCIk4dJ
djIydBDQDHnqpw5cVIiBE1xws9VBmWweZILVJWd4LMrx/g6UjyARrNPQlSFGZGx95RW+OpXxbumc
oqpLkkfzuplVoKGQLsNeMu7pv7p7JDE17R4/p8GzP92pXLtIIDOEqnsfTansHjMY8NfuOIPF5VFv
8EODAL3XAg8IqNNACD8Yy7mGUaL+ZnT8NJmxoT5K6lFZpTpTSHLYM1tVFBatbaoPgbCuDWyKgUIK
Ix6dsKll3+Lff12aNiT9dGQXzZRL1KHi0p9oXQXKceoAzi5unqDBP0UygDRm7HOnknpr0JKPE2tk
u2LNaqgarsBb2HxnnUIXBkxs7o6PWPZ/vEafYwMZHEyZR7yoFVt9N+kk2UM2U+pC8JaklgxFcXn8
+pq0dCG87cWgc3pPMhE55Jb47pn9Ckx2PcAC7KErRlTrYGyehpMcS2k9eJkQ1V9b89xOsm7unVAX
t7PtPEKoVXL4Ab6xfUOldW1Hy+nkwNo5RqaCTzDaT9FbijJXmsyl6cJKUAOv4INmfRKekhSQutSZ
RB9NSNjQT96ekAdu9pFECHhPbdMQyWX6rgoUKDxBbaZQ1PZLOpCikAjG1k481S8ionydesXRPVaA
wiVpczT59ocFASYTJRI0hpymvcoD+QPhfEf1/bphYIQUAiazBYFV0IFg5KeQCW3X+6ZLO+5H802C
/ldZSffxz+WY2KIwQl9Ko6Pm/LurxAawdCK26ZWAnsnZYEHV8XY6ks1sDozwaH0GkOc+Cvpo/vyX
NewU5i7WtKA50jTsqFGAziKa97n7qvmvUgqndxhbnmEJ0varmb2mf53tSpxNv4qcMe/BnICbI/qi
LhvLlwKjWgcohzkuN7eTlaCz63+wDk1hewYgXrWA5dB5YE+8aY6Mv2HiKvWhDTQZwH9YqlkL1kXq
wOlJE7l38/vuf4iFkyPSyQNp0e3TnJdVdJZ6CMf4NDx27ZFnoK/wCe/buNUHNhHuNbD7GTT7IUvK
oYmmcU5OOhWOL20SrLJsGGmpnGpcc9eAB5Warzr/kvEZLufLS4B2PaPgiDfaGd1sdPMWx8WWBs8I
PRSwrd8swGuxwrUEMxXWn0W3BcNearVBE4ZY+mosMv8E98Orcam/FPwSFe4wmemL/NB5KBiBHP7p
ibZHOR1dPaCPmw+luqwOZZoZEL42qb2Lpvln5Q2H75zv1prXOfcWQWwNAAr/f+1awa8dYz0hymlE
9igf4CWUU1QeN37f4x7mtu1LctsKMwBE+by8/bRLnKU5G8X5Fut6+xVegEW9e0GOK/GMmyiO73ly
OQEP9YqoNZaL6eQBvJ7ulo3JUTQvD++UefC40qWLZZ+XtZ7zv3xl5l5aGDXGcMw8KeY5Hx+NWYC/
ZWIUGSQ0KL+S9uBGgDhgFn111WSvTYJa1lnnFSWpkRgLUTXOhvbu7mdyv6wduf7Idhff+3PTC+d2
U+MiZJS96jGAry3ZYWd87Ol8pflFWvz6w1S2VylYwmc3jXWH4f1tp51EE6MlK5ps2SByLo2TOCJT
59SGz9zf1tZIWdCBQ43WMHzHdAnWa8Rd8zPCXtBxZhv2MFZRxeBMgbZPAkHPE92KbgbnqeWblC2+
MUWge3yzwnpzjFYFNDiVy77zpQItRQZFaYd7s+6NnZwAZpSY/HpO+kuGPk12VbxUaRTeuJfH5sbG
nhf1rBeNcXCCA8DQyPv+z2yHB/MQaXW8WOwA9OBxzIB+09HARx3MQaeh95IlRXLDVxCi2y77oAfE
RS33n6ePP1WQAvCbLcJw1tStUBkeolCHOSSOYMfn9tIKTluJwFdOCo9fj8vXmnB8X9Vwrb+qxOCr
wigNOhgeuG0dOVpEqp/oYdX1EYtxiVvweuSNxSNuQImH1rswvT3Z1edW795yNOoBB5UEXZ/s/2ob
kz7UYYjCEyZx5Yhvf1qED0L5uopyiCxjyBsFu8VBA1DbdlZgOacvaZcmd2eGMVo2t/j42xtriWx8
4iZ/ET+ZTfSK6BqTuPxqEdL8n/qLF8Q4ibSQy3V+LT74z19e6GJNFlBYc8iaymRi+ekYfQh9IY2E
8OOibgICKUzG5Huyh8D4UfKiwyn37ExJ6tmWbl0LE3oWt+X3oBYwNkCPmJ9VOcyWeWhujTmUPgs0
5vkQmSbfXIwhyJ5gY4SxPWjP4xj0U6c2KPlS3P26IlAHT2rdwmZozxuHzaJeRNMCV7xdf+Ahgzms
uMcCz/LEWn1DAXjT1HckHoTAc0DVkVgF59p/sgWblZpglMw6JHfup6k0eci8F334xTuXgcs94nZN
BXxjUzeQVKvOKqv/+Bp3jvHIMqw2NNPZS7m0jxZ/oFdSG5S8r8H7+FWF/bIh959kp14f8knoEGO1
bnS6m2xAnneDuZ17VG+ewfmvdTNXi3EpqjUmgIyd/b9H81xeCCJiYIue3ACKpyqJ/qPudghQWfZn
nykk0Szpjxezi2/zyGlPaIJUFvxlixAX+wtNbfqV3Y9tKFMXb+T4PZ7tExsFcMLMCpZYvCoHvc4u
ifcBXBb/9HhcC6/6jZ63axu2HrlCJUhfALGyzLYevSphQn/A9uqxJE/MKc6128FXcbjdEb6rnld+
YKqQPo1cvBSWVwVrtYuMoHKUfCrWBJ/beULRZ7Uq7neSbhFf4Ez2Xj0AFtsE/c/iPIGmg/NuEDw+
C3b1+Emxq/8oArZwPHJm2Y1YEsAYeMKu7nF/lCBJ7fZmSz6cr5zLEUBlUiGUcUarpQYn+TJ5KqVo
IEPziZtFZq+CtFJe4R7ZmpWa3hctXgSzNIv9x2q6ZxCu4uYNdUu9AYnHDhUVAvmHPfkPsQl6cgnq
VHLVtHAIR5wpMccL7cRvW5sZNf8PK8jJ26dKKOzbSxvbE1QkTeP2uGqRQ10nhQs7E4kEEhgptnLS
P1hWMmII4ZS7mQWUGvg1AzSKPmcWEYa1vigw9gQDUUSxJ/zaOTLaon4dVpMDrHqjsekN3q2V8e3S
3T79k7cNalVByaiTeEElVmNaKGhxGI/1uiWjjcJugm+9fyeMaizo55fE5aYLLyMRmFemy8MpINsK
RWDdZBkdZet497K0sn/fPRnFakNyqfLrV5A0AAY4pZVJ5dphYuPYz52obaFTqZ809wETLuXepDts
umazkIMGQRP8xS8Z7jt0V6xNNY76f/n/1oHc0Sm/OUEJcYbZLZViL0Oj0oWZUZ4gHs76gWznTE/0
4Svgpl8Q7IJ7bcW6Q+ZMIcQWpVED+zFcGRJMy3fxo4dPLjPxHCBcSgBawClgpzvk6LMcspFX/PZu
pd2YAiuwJ+ebSh/jVqKQ7XzKTU/Ve7bn8xxZip6Vj1Xb/UrIDGAt3L5v0usO/M4U58x6YfqOLUZU
7sgqNG3yjiRrDc49ZEHXEkxFQ9HMM7LLkTfnKBxhZSyd12nse70tUlKA98XFiNinAKiv1uFtXFBe
lmTTab1Fi9xhh8BYgpLgB4rTpavDBxmu8yjWu1RZu4wNiK8xXinrHU3sr1exmTOAKukIyM4pIflG
+C9QCoOGFVGJiD15d2wn1CyrOWWWgX331QDxJPGQcvcoa2quSCTRlX95OFLtfmqaTuSUK54CzwI3
zFrzrKzCvJ1tp3V+T859mEtjJeR0JASgHRs/yBYoNJ8qtYBVaIvzL2GGb4D/o47btclVHayuhJEx
558uJuhMHDP/lxyKTyldPVcIIxwoIFcBZQnW4zdNhyZxxtkFROr/9j1umt71Q6hLlyRaQC86QJBc
pmehiTfXlZ9OuN/clqYkmhlDZkJC5DV2lXL/x7Ce1tSeTYUU+5GRy7xXCCG5uuT5p605uzI7x222
GDMbIOZ0/iVop1zMZsBz9ZQP1PRZm9U2+ONFmFf6Bxh9G/loXBbA6lbD1JOFkbcz9FMIA0RyHAwx
soaIl6kyEMPHdZUBySIeS5pwsg5NHUssIixLf+J9dnJYS2fC6mS3bAI9JAKV1kYqxVKvSs+ELYlT
ASEGwe35yivuYrhQuLQOLvyYc6K00+ngk56/8zjZVvKvQ0Hc03DlWFluRlgBHVua4nndYsdgHZJP
vV2ZkWcW0U5UTshYXLirx5IWoR3v1PtsHsg2dxQIEwZluZjg7aMK0XMVQJ2NV61u8aRQfHLr2V7U
BCWXWKhpti0p37XlypLwiPatIVYddy8jkWz4cIE9ePAqjfqSQdyiXeP0xwfrve9y29nnNprv1JU+
kcff13HMH7o5sL+xTKoUr14TXChE1vw89++eh8LrIRvUCCQDrMoZhsRfJDWuIpPj1e2J/tM1qNo8
dYiuwjIgG5M3GxcBKE64JfGIL+v8sKP2lTC8frz23JJP3+uruWNiD6fQmRWco4v6fdnTWv/gNc1/
qI9r8Dukf8Q+oUI23J5AKjblCSsjjd9/tatipGi8QbOVI48TdhuG2PbE/dOHQTsH1zgKMkBTuayh
smmTbskwxX57oIE9PvrriJyqlroFBsOTsJV6Am2Sly9osdlLIO6MmkaUPDqDLY4ZfYOae9JdwJaO
D/L/bRP332XhbFbzZfIhuAUfpT1tGLq1JFXbpx8UBSf60e/kizx4iW6DfL2bxJ9FMpQ6azgY+W0Q
oHBBw0mZNJlwvP5UeIIZgCmarIvQm+jsC0gBjktndDcQwOI4IUsl5dPyfrHEohfz6ZBzIsPfMYUL
GUo/qmTdJKOGPeLwMdn+AHyRhnuUhVv4U0KIpOtoWkfUs07zLKa4xVs1x5HQ4i/9TJtK5qPGp5/y
6IBGxYVoT3IHThb5Ky+KYleYqS8wdlWscUcyRfov5vE781c4p/sCrFLTzHIMVL2VFeLYgtPVMYhj
0GzqeuLL7uSk1NDwJJ0lQzsbXq8TcziWlBVuHxcsUJ5AQozRpn8FFXn9PtQ59FFVQnWpE7syumdS
ivAW8HVEC6kfggRhEhIXGqToqLT7+1kfrguzJGcgaXWt4WPsLve4lQsFns4kChl/gVNEUd0SRnpU
Oyhr/tOBQ9jnGqxwApdndHxGooJBDc3jtobjKVgHxCeiDrwThRt2xyXhLxsSE85SXu+VHYKUmahz
cg4c08ToXTSgkFkcwRsocdIkVfYZuvhWsqI1n1Z9+euF5HifaE3Ct0T5KHrATHpWcBpXtjj9lDW5
hkqAxdtZiovplmTLOtCEnFwP4nxugK8j58SDYsrfgVFXAZglFcyCdUCzzK0ZxKzHYTivF3w1RbwJ
kS8MSkJuwsUkKhjd5UFJfMIwyzg5Oz/5KfnSaj2a8TIgigcrJVSZIOSOBlcWmkOmwfdd9jEPRqqy
V7hzwdKCW2sTrvcF47HV/xGi1WiJMQGt1NgIOZl4BOK49f4iLipLRV68y14oFIfYQ+iL+8L455ma
cxbmSEsPcdhmTqQuYhoy4k9Pdh7MP1e9N/yFCEGwj/BxWN3HUsn7cXgxBnB7mhvNtQeM7XaL/baT
DCLJ++79AfNCV3A8ixB3nhDzS3GDr7rg1aOYkGuToc2i3nCar3GBbht3EM7ySDqlCo4obvOtoxIY
1xPghNOT846/DNIrnaaMG7U/zRhYibBMpmZFRGI4AHCpCyMZDSzZNtDfwR4xLlxQffa+G/EueKdv
9adHhKP729/ky716F9x7xnXFmm2ct/31Pg9iPSer4ul621GAQsYSHdGqbEEOrZvikuXZuKNgwXt7
SJ4V4WfHtwg2rCa8i9J8oNUoA9ZdCxxAjWUbdFwYmRZ3JgqAAdZMXYxi5yYzxwYfcdoDAbW4H3AY
TXh8aMTBerqxoVEftsT5UOJMqO2OJVMQlmcXNrUGb544jd0QPgsw6RvI5073kcSo7HmiN9EQmBZV
pL99EwQU1KYfwFJRCVmRQHJlVZdr7iCfZELlFLzHz+XqeQe371h0ADy9Q3+mnKFy+zmunP8P1OxW
12HhJdMsme+973MykA+dlGGL1FC0O1yZHwushFiHrZDbHmRIV2oJfTGGQoyhJWq4lvmUGNESSn/M
XQps0PmGnJx5svYZk8nntqHIB4CQMDJXICleDPMMCHGUZjcVVBxLzEXXtwTNuBhGCCEViZ60Yimv
xvZFj3eDScrOfobphdgcfj8zFXQdjjYWHjQ/aOEXKRzLUAdTmFCU04LjsO/2BXeVBPXPRbfa+TUR
qiDrYtzrvt2Lp5pQXrld60o9BdHXfQUW514mzenirF+lBgGtmeWpzCqpmw5lkbn2ztnyU6V5UFqT
9OKGH+L91+n/oN8o6S31Dj5LO93kyyNivAem5U8D6RIF54AGb5bET4k0uDHgvc11Etm1MdF+0uO7
G77aD5BsF9ZgcwpWrE15kzwANpH9TsU2oSXB5yZwyA9axrvI2Iu/Nt0kX64I7afMlrLtS0vwj9gC
hssINJL9qDyb7HEGjVdUSnr+jatKQC40FzoqCIurzcSGC+XrIQh2d5+goYDtUPYBfQMpioiurGiJ
8NsRUjQzhQf7D9OuP/QTRuJUsSWBLtfR0W+3iLwkTFKc+Mos2REil2aODAHr2iNfgh5LPEu8LAtd
t9Mowmfxp6rG0jkoQJZH06HXa92Uose86YheAEhzBGuEBipk3kBhV4MZY6qGKiy4S10X/Fo+KRDL
eJoQyqNb2KYUHeBcaFROLOTFX7vPMO36wKmmiIwuVjbrFpeVLlcgMZhEKji+I0dVNeuQVeIBxUCS
1CR5Kq/gHeTvYXQnK2p3ugy346Pb35tIFd4q7KeX7z31Wz8bksd0eVObsHMRWaKTG29u1pEhGjzc
xAqAON2MszmaEy0jrQHSgupVA+WkozPVHw34BSgl794DCoTkoJ6517j3li1lanwbgbClpxuVtLhG
uIh2Lmi8WMbC3Hn+M9040Axal/pQN5AjYO4PbFTGk3/bGoonsbFqfkDRTnhH6pYoYM9iqaevfk17
JX/VJmn8sQJSOVbtuRUMybrbVI1nJ9TiRI1ChKFHt4Qy90g+VoWkJ570IQwOTM8aIkYd+lcKeCG5
2atmcGR6a1EwDxub1DYXGQc9mzze9RzP+gvqPDu8Pl9VEEiHSgNnr7qRcStXsVqOcq8fc0RH1gN8
GpG3lPvmnh4GY9k7xKPPXcw+wBhfy05njCIoNd4VoJZh7oIkvEOCcJg9L88LzYbaWvLVTgPYuqwz
5AeKSB/4tHfx6TLx14kuWdr5ZaXBvxFuuC36Ny25WG+dvEzSN08bUSgV0KM5akbgZsZShxZYl+X8
8cV5Eb3ibeqPU1mmloIE0k3+IsxGAfy18RUzAsFFyEY9ZVCBF2HkIadlZdSdXC4ahssM/vPqlzKb
qKHYUVCafVo0f5j1Y2A0VcV8gBr3CxNy2gCRG4FLxlxERZVF/W6q7uUOUl/VKUZ/dJ+tlKE4xsVj
+UWK9OXF1tB5kte8S4f7Tt302tWJFZcLLnMZRYdTnQidoiq0Vw+ZM21zk5KLcplr9rmfOrmHi6Ec
kPx7ulZshEpygwudKdpIyoSRGGLvE7PThJUHI0XrU1izaAP87kcNpiEw+NSb4q3QHeh2XpAqE4Z4
Wj78bL85vrTbymQNX8SMbCUFc5jtZeihu9RYzwvOfw1FmFKjpGHxjVgOrG4/OArC916q2NE/qTC0
DJYK1HmsI/lQAaPpLrWA+3e3evUDU5K/VJL1nF33rvKtPrHRd5QQcrWPcdmlLWii0sVH8kzyX86v
qAi2Oxxgtg9ngzs31iX60aHIpzsLUOMQWCv1jep7UBTXHoxX8UqkeTrM+HOM119lzsy2o46am7dL
NL2jF/dvdHTrpXWbVnqoMRYztQVVuj6wtuLaRBAO4wNyMB0N/MfFrvkW30JNBnSksmOOfsbOCPUT
Lt4rxZxqsLaRGVgGflhI464z1chaAngfTsWr325tyVHIs1DdmcSJW+B4JZVlQFxIu+7IGETHViLH
RWU8b+3u1QKlN/tl7wULoU50HJDtVmKlLVjcjMMPbk9NSKNNPDAzdnXuoKa45phiwVHnlzTpd4Dw
0bgoDhGnMwACILJkaq/Ed1TeDKOOPcjpN7SgQYAES7tRDtyOpVCtNcZJv5+LOfRu/rPYy6+R1c7o
x1uCiY5NtxoCGR48HbvSfHccK7UGnweLhp1KiW6T8sjnrQWjzwNRclK2n9uIlMeqCY/v9MHCfErt
AwtLEVRyGlYp0GBEja740bs4i3EtOvHRuCGUDEasVnQrE/npEQWPjVz7kWcCNS5Re70EE5q6khkA
Ce9APWtutHbRcW6F51jLXjqvj4Q+QhF7kt5bxHpbZCaR1tbBPOk443MpKDahroK72cH6bA2CIm1R
tsp5h9tF680eqz6h2B5pF0MxecQE1N+EFjXyp/qlRlH8YvcpxWG+nS1reOUK/3yhkANff7aVQaYl
GP5kJFJ10rok/p5FLuF74/ldDHd6wQ7DkKR+6+mhMyaEJJnfwHlkjjyjamRjmMbUq9EofdPc+Svv
ocpgrTy+IEdOEPkxsLF47hJ5vrffHfxHP8yiNDuShCeHCyF6W//7QPtCSLdtudX2HY27ldX4pomW
QDrPZdE9+UazzA7Q89ubcmIVPah40q1dIMt4/tGQvAk0nFZrpnn8yF02g60paRC2tAHjEXKMIrDQ
YC9r4Yi748sy+OqUznqfKEgp0jMyjxKwukhY1Pid5LVxHy9bAHqZ4W/aDe8ThhLJv0jiG4HD+pNj
c2Rlfi3fHYyr656yp8jyS5pawmPLbI2knCkZC0GhNfT+UXWvdochciZDslm61D3oX4c2IVJbMtd+
BhKAaARHT3cK6EfPQ6qakxo0xIIUjRi+BODAynrMTubhPfkYlqaGXjObTEw9cYNZxzUwfuJ1pPyv
mTYu7TvbwVqJtM2thD1qj7B1rfmMl9IJ76j5O3o5k/triL3B8h5zjft7Y2rqUWij9ey7x2wOODqE
Lp05XTLVuk7Nr6reVtMBystFk1fY8wcO8jfRS5mVOeQaMXMRtTGnhLuJj7e9aalfsOJYduPF3sMQ
1q/cMQdsJh6UXht1KfDEmlkp97YmfGYp5ssjacAw1i467NiUDNkPEpjkpFVo76XfkgeRGtqbWwST
BY1g9XE/PxzUwbaL5JCJlP1BfWv4VdZm6JEfjjBJ/j3OZmllEovZyBpmhLAlkBzNrgmMbOIgvVo2
wI+XyoezeWCbd2KcJqGf/JGHlST2r+2SWS+Xb4tLdamBXUhAzfMn0bbSH6mhlL1mdnkzGdWEUshB
npidLZCCgiHZeV7zGyp1G3ur0lPk19aVHpGkzgxWZIvfEQEJT98DDPW0j+6ltu0kW3IURQOs3eg8
DCyyznJLOaPvwcyoKPbYgHTXFMDD8rbq7Dm8HIYiI+T5wCiJ6b3a2IYjCeOBqgYAPKe8X4kXKTdm
VhaN7L5IaAtirubEeaTpl4DDHN52ldUI8QS/V93/eBccZjRqtJ9wwHrlG7+mutKZL8O/uSvQec1o
EbE5uAhk32onIYJYMHfGoCtOjyAwnf/ObEB8LIB/fOkQhhCXpPMqqmeWMTYWSPM3S4Nlm3Uy6YV7
KIaB1geySj/QfEJ2fkX2fpxp6ER6AS1vdVttfw0y3RzWBZvbhjEQVN1NCo8skRGRn+c5AOjDHJXa
eUlr/7c21RVQVJHxsYoP6o2OFJMho7jb1bLLKySClvqI7UqM82ct4uluUQ6uESaM08wQFAsDyI/J
aFTwGkOHnN4pU+9yLsZ3qY4rqDmmBlaHxinx2U/LOvCielntZHv6ZXOFUs2X508HXs26qVCLDDuw
Bw9FVhHz+CgSxCUqRXbuXWHRb75ePJhWHF9bwqJz+nZ1iP1YOasLfdWKuCZX/dgw7vxB520xtVc6
/6NTm7AlAXYTsu1lZdRv9tWhF/MeGTrqz6Ln4mpyA6NQPAWOkWBzJy/dURDT2DrMkyAGchYVnd9H
dBB4JDnqjsrzgtfGVf/+ZyWDJN8DaHFaYe4AhTYyvPcxpT6imOfePxb4GId2rzMElCgIYjdwul9u
j9ptaKGKH0hM65viEW1bD5SHdIBKAjJUBMjk1lQ+JV2NR8SF01hg9ASFx80w3G4HgLml5w6w5Vde
tnlNoRt60i6llH1QK8MpX6ljhZ6JrztCah1wyhHYTUedK/udQ1kPq0m6jVztFdZXSiTfdsFDSOH8
tCdwjk4u9r1dop8pTsUg2f0/3SBv2RQOlFFYyFv2T1nUm/lTEmNIOymNkmsW0LN4h6B+quc/OMYG
kkwUfMjgRrGL83mxE0W3zRcXECvbOcMzQ0Mpf1d6B9fTxoD282Zw3XNZp/raghwzrCOQOH+a4GRe
o+yNmrKvv9r/Wye9FAorfo4X5OI5QMX8jM+Dlqz9MJeDCJhq27XFQWkEuV7GjPrv17Xy3puU7T/K
lWjiFblPRPmDnYLwkOEg3TQmmSt2h6UzHMSsoGHXTHer9w5vRi5o/jzsGN8LbMyLJz45s+tzbN6Z
/lD54PirKy4WlUaGtfAklF2SY6atfG1Vc33R7chly2PFM4XyP5RAgCA8wxyPYITfGBeZ/xAqe1ym
+lE3H1Q2rLaLs4A5j7fJ4k5FUEUfOHJOkDqMaIEPjyIH9Bo/W/Kp6/F1Eh7hDS1FXomS8vKPO3ql
N0dugWKcg56pGds21ocJCixjWCgun0GRmllSe8fm4mMwrik23krskCFE+v8rk5Gu/Dzq+YDLY2GM
yYekcIb6f8UUKQger1mnura+zLRrZmLtLmt3c1L6e+8UXSw7x+a/0zub7z29CeWEA1+WVhxgPO9K
+4DPEgy4VJGUiIGRDlHKmoGL8vYardeKB1YrDPP7lpg06reTxubdZclZkqL43wcVy2Y6NhhXfT36
k5QMwsLzr7YIJ2UPOwzdZoe1mYtYC7U9QUb790ZgiJzXOH6UsQZiqiIf3ApVsio4aWV+SbOTPutm
EcXX/euwMK7h+seIbVfbR0uwsJTulTKDQALD+YPshfJ1HowreCQVnKDWXh3IEHUXc5tdXscMvMmm
wDPyA2PgdgoN7eImOiS5uwVUMdyAyg4be9RM7k80pzUwekvu6p4P0HWbTfO8T63b59KjZ4Kltugk
NbAZF7ulGT0cgKtVr0sOXgF4NpFahrJe+fFpW32LYL6n+XNeHbPCNqEgTsDLwxPFD0B6SLXXU6Fi
7sJtUAigjkYKqf9TPiuEWzDHIC/MYlSKIz4rsAmAKt7iFFIiSwqKbpNhRMxu+T1I/4gzoEX+T6Tg
M2LsUDaC50MZIrTmZxr89s1uEpdei48z/yTYJV5kmg50HuwldjJ+awL6nHZO/yalUhe2zI5KCnxr
KvPZzk2xGRN+FsxaBCZWM7h8dmNswZYBSRGi0AeNv8nDXu4bAwSPYfO+DqckR796ftiEZI5UhNxa
gVNvfTIGhqg/nmsaHt0NlaokMTDTH2xIOXeAO5W7xnmxrUZQp/dIQToaUcS7y7dg99l/qx19vmNy
ei9LBTPg83XVZn+yGFyjd46qd9qHIWhjszfuWBK5fzLsgeF1mq7EHz4XGogBkI5H3RqCdu+GGuw4
sBScVQd2UQumxD0bcgHPufMtNXCMokXs4XMNtCB1f08UhAOpEBsxXqlixFvsUGjKT1zDlFYsu7xX
IDhkISZPN8ZFYz90dd8/mEMTG7ruwcGTqa5c03JdsDxmOimBhf3c180G51UuMjIjKT5r3CJ6IWT/
ZdouTV/p8Q3NvHsiCkz7px6zmxDdLvesjb5mMauszq7EIzquvCDT2FUieXkWeD7d10U3uRDmWScJ
nYTiTpHAmcnne3wzxn9m1AJ+y3bxJNgeMt+DJZGcidjcLnodw55OlnV+ZtVMwy3eUuTvEK6+bkOF
zfYjNrTTfNAlmHzPn++ARI8U+NcjJnWvhYoqs/G9mwb7CjXhA0ObeWkre0/0Ps8MM1OjfHTaX4pI
ZxC6FM4e5huM606x09Lvb8GtzxHM8toParJeqzh/MXe0WQLoeorWafOcbAkw3/DK0MEmIG2ff2Zh
8SVXW64gEjiqsm9k8dRxhCRbRlCXpPJVCBzupBAN/jQ0C7IgptdQyocz5ba1zg6LvwTEJS2Kcf1J
bQNZAxwyosWQGoJ86IKb1k7RUSfTwgeNqmieb6OzW7CUhukmOfSmx77ECHkMSyEuPs54wBP+VYT9
Ol5S+1ADjPQU+qutNtcUloz4BT1PulNOc+eKAnFNNtngm73+GBehkrEV7OzdMoypy4dZtOk7jYBW
tHIoIG89wdoqwnBeRuzNK5T39rs/iRaKB+cn4/3nALM8EVa/RkWWEWJY73ebxrWbSvs0jS69cSO5
g1GqoYWxAuiIEmnQ42+LLcJuskNcWQptXofqCWdgjHizWvwj7xmn+yG7XcINuiGWeQa/PWQb8bj8
9/zhHELUZVgrcY3Lal33CMa1kHVGduBnGaub4BRWqGZNB9TecVm3pcc4lw+rf9NFvH1ZmIyJCx59
t/VUiraE+nvVWUHQFFBxTXVntNsBcHO9T/7N3pJ92s1V1kXU5SrPzaXnbn5MvCJa6I/DP2f0YNUS
1mbTeDHFx6cETKeZhSIykxDCaeiqSuX1YA6v2b28VgjNMUM119Tmk88w8pVQeeCeFh+0gbFSkRsK
DhvYwBFFDhBBGRx76UIqOvFjEIDOydnRAXA2m/RuGo3QP4ScebiaSBXSgCcgCzxGXWQZT6EJN6T9
LTTFG4A6nr2tA+udD/NAKo9nR/hpdkUD0ql8hIJ3bp2OpcIFxSizfz6lqoJxCQtBD24Lidj9j89Z
M/iTrEwd6g37Og478o07aoOXsHtYz3hg894DuuAUt2ZPGeQCwfDHjKdKT6wa79+Z01cWNueV/O6q
L0Pwih9MSGtWIAH4smIJ/W9Lls/53eEq7929C/5Fvev5H38KSYCN6vfDwe9gAcBEiDt+iewRiOM8
n3GWswiTFt1NMIVLcf+NHO4rJuySUKXkdnBUVShXcGLJ+RjVfDtnX8RrdWxqsvfg7+SRLjX0gI/8
S1dMTzdaQXw1YirQkKfX+kQM+CUEpNtYLthOBpDmyUBYQCKJZrSsWEcGzb9H5PokJkEZRcA2/GT0
DoE3yiJ3FORstzhzpifZiwu9d+tLLzIu/DijASMNdRCTrhZpp7U+Vonzq2ZyWn6PIIqSg5qpdvb4
cXunJzBdXXHL7ejWK/yH+YeH2RTQn99AkdlfkHunsLuhlWl5GY0aLYFE/x4OVKdpksb8Pas89wjk
eeZsUVS3iHqm30RuQmn3WP7jya84p8uLnojJJhYVqtnZwcfq/bT2cT8dUFOTZtp59qZmEz7Llfrf
sb1WAm9soiIJrZHuU32fyMYxtgzINttpboyJrt9xIbLJdwt7TxpZSAHIRJUKzzZeV2GXP3MnWdqs
9K9zv3M40FXfwkdOw2N64tRe3u4IEqg7K/M7TSPWB4LoNmfBlNjta4rm7Z1C8K7gd1f4jupfGNea
VQvJHbhaTQXWcXFIsPANVUOUDuB2IhWzuxHYwQdaaTPKRCA08eOjY/1MgTbJcvHaliMaHUPBFDJy
kejlZuxQGzttb8b5G29sNpNn0azqSbZIWnqu7wO5Egwv9QAXv3JBxGMcVWl7GruI8iabkDMPcf2f
gsdb1edHFF1/9dTwLZ5pKYM6+197rWEFI+vpeszPVVkW7QptEFstrOOvf4PI44yJWHp8tPhED7h2
+OZGqD9S1ebGRpSQK3kBdbrz887PkjGmDM4v+XJfNIb4y/1RVsh0J9H6HQCRxuo3eDk/f8tBLOa6
3T4py+50hBhQd8XqR/mA5NwJ3lNDGSHdlU0mOg7yOjhN5HEpFu4yH4berVi+NIhUiAzCjTiJq2Pi
Iv7Kb+BsWm91mtiQxqVKzbyu9LKHpNJigzZ5W+YqmwZPuL5qt0+0zTQCc7GQf0Q7bxUI0apZv7Km
pj8Wt3MQHAz67hwaQbdAhsBHziQ351WeFjSx3ZCANPYECexqreMYJhxFI1+6kOtUxiKuDSuNrEeL
YxdwpBJf9wnsn1w/q4mny4H/dLhF3lk/uJJh1LAAovtdJ/fo4LVZSiIWzPO9+QxFrgnzoudcROua
EgEhXc1yvr5uFJNIXCk4ZzBxOqfH8QxnfAIi0XeDmHXu1NRMkBSqBe+rPJ03gQaySe1vzZf+vzXl
2tp2K55dAasNpPDL89FUmTeOwqeHYWbHHcxcgy3d85fX7+iNwod5RDhLlCW4hS1/CfJ3myA2WvB4
umW4n1yd6pKoYvwF1KMdr/v6LOsRl3rPvoZWlbh8okuCx3KxYEFdCZrZcOcPK2kBwBlK7vos5Szm
39lxnIyTx6z9HJ40V0p9aldB1eUO73/5hF9uHG/sZlXLYEva4BQ0pot68bbC20Hs/GNpq+u8jcXD
P7dWj6WM8py9Mt+mEePHccBJ7vAZRCHd7c4arkJKWVMdAwQULVMTLc2X6rp1Q8ym4hITUvJD0sH8
LK3LJT0bD/hJ8ALksznLwF1xmU9RbhEVRnf2VecpciljTH+hEn4g7hjKqMIlQWyLdNXKiwWVSyPx
RXUWWFHwCt3X3SrjT5pF73oxG4q4dB+GQ90FLSTCEqhlREKJp5M8fjK+l2zuqm03ZXrSnsiYVU66
z1jU7Q35zx1G4KsXtV+zU6T+qvXoZw7XmK4/SLGZsKo+jWN9sU/U7CXdHbfP+NL8KZ+DHr1IC6c8
+U1oD6Bix0kEzK82K/KVs8psoqSXE+6KysL6a9TxHJ8JT51TSynQjpISl9MbxfhPtUlSSIAa6roW
tbjkjcMTHmD1Fqeseti5dfZ3vwW/0JFLYxD7b6cvSkKMb4lAp/4EOFafiHAOaYJFbdlhbS34UtIL
s3W52FIclvlxSqU34NSk8SGn/f+CNxf6lCla+MyjYDRQfDbVSrWgy//Pei7MxHrFoieWAWEWykLH
AWzxQSZXWh83R/za5i2bVDRk7VHz7/4WeT0L8cCirPkGTUVccgL5bMcPtI9SHITHikoZ2hxpZ8ML
l4jJbeycwcPvsTPXL5vjC6rpRHAlJj5U+C5ztiun2/DsG9MSWgLqaZ9IpzWoAFx+73kXtL5RTPZ6
HR5xw0DFABSuoUxLOO3o/uJLsNCJRh4ND3dI6rAlqnt6ZtVt7OOvBDHGVSAuU1wXrzWZ+IBE0CPL
AQyUCXtYZUD/rTqCDUSv7DoMk3zmas4lyGBUeLi8ae2SZGnkrKIuKOKJavcDR4iw+qG0AlhuEnS9
ORDGmZYyK5y6Z6YCyB8WknUNxajUses9WgN0H2DxtmtrCsn9794L1UWpyRW77XFjtWVfWKlLmheH
epoWONSXiKlYXo9uHQTiN9XPT+mnmqzH3ccmy+fyOpuWvPCHihEH84BYg4vYgoutT7QiUVIcBNnP
TZSWqBgnJpx11XVoy8QVxzqmiaxny56qOPdNIALxSodiPB2QniKm3MTxA8WMxama9d5bA6E1ZUhR
qwRm/mhvFmSem4UG76nfu+1WClRhCGd94srRSVVaEsVPZP4CNlO5ziZSlBgvnmUruSbJo97Wxued
+jASbFt/lbx366hAwxtpiKj0dRTuA8mKoLyO/TEm/+CNwdVbMbmLNokfUs0qEaNbKU5xP/pv59VC
o4Dk3iDTQW0JfvDtjPKPZVcX3b04bnGBXpOB0AWMCpjJZ4CtS0yvVsdpx9YdVE+rK4h/Q8VpfKLs
OoS8GBx7X57P84TVCXtsQwiSaVgp9smW9OoNmGgyEiyEvx5Ya0jLjXN76YabqihWvBVBvfNLdZXE
szXaIM+Gr9mgiLSepfr3lQqdMBLdWe4ZWPMs6KAP3x/XpVvDzuEWcloF5gEUixHlDN/wAukzlDBW
6bxc5EbEKbcYRK3S9dPkL7o9Jzsmg7H49agHbBSzsOGDgO40k75BpNf8Uvs4fhYomxsXVxUokfCp
Rh6sLci/48UqdWvooUlPiIi55qb3VJE8YJT4kYj1CGgllSaLfkQRn/+2Am+M7KDw0dLvsGMo5NjB
+1AgK+xSdnM0ympyyCRQuHxnupLFTRWGlxXh4ceiNg8RLB8iUqozQoQZgiWeYYmS8wDngqONt4Zw
0U2JDknLndQC/1KJ0Ft/REH8yuAUd3i34jI6+B3YQ5QKFEos5DHZFParHzBTtDct3vDa453yhfzh
FQzOxMmCVpb8K4FWSBG7bqrnYqXfOikxFWz/7JfG6Y9ILLHen5KHE6oDaZRv21DJetJQM/7lPM0W
8zfOStZLa1m044s7FMVoZjzcoagRkjCfNwJT+ZYwaulHCPjOUobcgMCKsCmEmIccBMVbALFbr5BR
DuDebjOXmJrwY6yypCfVNMzXeQarNG9uxZD0Dpjgkjyd5xLKWLu/114hBvt6NmxYfTLMbHTUFa2o
VqiudxvO/2w4afsjwom0DPgXFw4EOOUlmiw8Nzg2CvXukpQI/UCX/5LWgIH3aSUAUUo9o/JFi/3W
7VgEW8WcDBOPdqqdvVg2bWZh6rwwbWwncUz52ZlD1/AX815Fvxn1JHb8GDePBARw4ARDacwvnPIr
tCRHvEPxyDQSSzkMJbNEWbPpAlegdPZpWO1lbfWA0PHIDkRhImf9ARuIsrdA6a0GvWGn0wXjc2+a
gsZmSkDwW6lv3yKZ74zu+pb/HhWfNkzk0E0LoqOH0HbLioT+2buogPwqMEabysxbTpg/jDhR3amI
qJekebybgWGFdsStGpyuVkXnFpXKTXs1CmT7pn4mp5cd+gMUHqRv17+P8N3NyI+pyndmAr06rAVi
XKapKsLafdyj0u3JHSXgO4vu2a2DP53AZR4nXJTNqkjq8JLnMFGGz2n4fCAF1U9clhaxcl6ZRoQD
dqbI7+S0CPqOqlr/J9SXZmBP4YlyAGKmIHkM8SFB5ztAkGRlVRN174C9kbkryTVN/TqEYl4D8EGT
Di5GhcKYw3KB3aA95bv0vgbfkiotnN1/wNruaNosl/NbTs0ZRMf+yS8d4Y7Z5+gvO5QzsK7zUEni
Rxm5MeT4Xb01LFELuYN8FlgXQ+WDUhQjaH8t7zWYLAiWoASRtZBFJbH3nY13t06zgFkvbhkbkpSm
a2tsin98LKurYZpb3pKnKVmLkRTcROhdX0y7L3RzX3ho/IN2uAsDhKLQ4ytt3+0d7bFIEttqXrlF
RmLXf0ALnC+rGU9e+3mrOB84qb1Gny7eD1NndJKPIZKLOZ1PNzDslTCt31De/F6RpDOv+5hywLo5
SZ+SzbWsU6i+sVIIUzEcb0A682GKTksyQsdftiiXBhGRCiH7BeuIUJ57khdniwZ9DkpbN7wv80tj
borVw6zIyOLsj2J5TvEDaJr8SgFPdR/tfaG4Pvy4d1ICBk2e+IH0jg4VqgEggnB4fKdtTdjQb7/b
lQlzJiFd8lKl8nFVL+XJFrf3ofF6lntQCcEm8/q5eLM1M3wt9EjFmeJgXfWX+yhjCstERS/ZBZOZ
mnhLMKfxjzVUIIJ9fd745G6MpreidBzNYHnCAMYW8rQzXrycv2iNWb1+XJoL+hV7eV1+oV8fbZZ7
eNgLuuQekgGRBBLrTPK7g3dB/Ubb340d8oo3KWEOvgim7cCNCoAFkmwMMQr6ONiH5Bvcawx1zi8Y
z8PRlrRpmUdHqFiLndzQIDjNkySvu9cUadqHFLpfVMjit2rgbLLFC/8C4WAGXEhMDU+vrcb5vAU+
PsqK8QO+VOgZsKzfAbI9hgAbA2o/Spd1fJkGuOOogGGyH/tMPp5w4uxd89xZXgiuuoqzThPLKPl5
Q63nMwznWWRz7QH/bF4jUfDZ0tNxdr6/AY6PPTtZpoPBWSHWSGHew5ECyYsI2yCCXhqQd4iI06HD
gJ6iEOheucgAh2SLPGGr/OywhlpuAcUDMItiSrrEwbDuq/S8KfcaaayF20ivwYl/NHKvdgWbT8CL
24+P+1XdtKqq3Zh8S0UET0U60CqWzoJB/RX1RFRFztjgAms6RBa/w4ZpqJ3yeDnn7l8Oynw5cFQd
bx0nuYKoERhIjU+7JI9ZtZJ5c3VFGQaxmCxgo1U6+C9wRG5abzT/Q0ZRT/55S1/Rt/Le7rAJLzBe
m7ExuM84wMQyx7F4D1iZPdONXYRJFFNVTGtwi77/4ufbNvFWgQTll1MMK5kUyrZRgbraFBpYsIag
8W55jayfFTRDCDaIB76LfDM2oFiaVu5awpyxTMXkMMIDwR8+kz4VjM0/hLliFR4GV8giC3IsvWl6
vaS/haD5qZ2xdDHgkxaOfZAvB7ESLw1Memqicj23rv5+kFZvSgeXGSbEQMxXI6lyoTSCA4FLy+N7
lKslr5ieKfFF94Y2GpdWGkfdmF6L//JEEsfKL/Eu72q6oqiEH6eRR8AZivnBoJjiGx5/96ZOL9r5
icj3jgIYAOmQ2YLmgq4upoRxOr6lkwVn5bxF4WN/0lzoDkUMGQxI0zzbydhLvSL7zNmsm7VB6nO4
lUk0e+9dUrApgtN+2h6WxamLpnqJpxPPdLVN8brj+LQ2Op/w8lGQEUzA2c5n51ybbj0Xk8F0nJy0
XN3Jw8e53rivlnNNIDuQgKTfOmF/2jfQKkrA6sMNkp2uOC3F5GmkvYFw37jPpqR3galjvEYwLKVZ
PZdTZz6f1qyzfaPjflduJzj1ShNB8AMB98xRSqu8A3whrv5yeMgUTeuh060WBDVk4E27e78fXrgj
/jx0+6JT3sBuwSXNYWnYhsQsr1Ip15xescANVFGlk6EUKih/Hlktnnfh8p48yl8fuiup7go6LQlb
uiLFM7kf22GTf38zE/UJSx6sEgryUg9BbdfbzfslhPn3beX9poV+p+CyEsg22y4OgoKW0s8YJGMV
vwyFMg3sabUfcsGwnW3VT0Ct4oA3Rx9xunTFTBzFinCR+odat/cVuhm/nOZfKVxYNcucIZMnDcwr
UgH4a1ib8XtpJ1EF/ObPJF4GA3oaByrnMsbkdxVRW5RJYdnIGCFLQ9m1Nit+lHn+N0a0iQYIfDbD
h0YkX1PdskQ725NMLJ8pdKceY3jgV/tksoJ9M+sEoo6EMbbrsyIfxOBh0+XLFG56NLEjH6kSYndy
I/6MPFWkWzB6A9Wu3NL7gfxfmeVUSaNKDCtNJpm6GhgD80aUbwOybmSWxnTJX8oTO/lnXvVGdOUK
tLQEe/X5WP7FNTMoy5y6b1iZjhLmXhDOKswGr4YsE0f+/oCOnPuW2E/q7cbJM3H0we41unG0mz4m
XfY4cETQqwIZa/sjIf+ux91MvUiIGlKlFxxzfjOc1nAjA/kKlh+yRHgShEadPLs27a74y19Nuj9C
ymro+GsIU5aOWh398dwfIP6tZ7eNwpSMgqnur0p4WawXkjvHUe3wMgi+SMZCk27kIeB1VTMAxL9d
1V9J7miCu/jelQoURit6CpVKaVQrlZ8MtkE2t9pbpfQVM5USoQ7g2wa4EqILTTQdNMBqkHFgDVLR
7DGso9iNEuHseGur4Go0F0h5/E545klZIkPHmYHt0Shd5VcnwtBVXjiZNrSvdt3dp2Mk2DhHbtku
aGeWyoG0qlt6qlLfbaqsWnAfPw3jXHZpAtUriQUuJXpVz++xQ7mIG5pSY181WYBYhi4NwREyJK31
8/fWz1i+taBQd1LR4ExFIObCCNtzZnmYKx0c1O66pMelsW97Q0spzL0gatmh2V7xugXEMn8JGhB5
1y/zIb/KMryPCQXSeDLZQgMT7gcI0Fqnwvukh/kbI8fAURfDg9J8+musx7+9UVF00WlQfIYC2bM0
5uqBvzmrUnNL+5RkEtLg17bEHLH2GD03nAvUBGO7wavP+QhysuEgHbIoxp0BG3UIineVBlDkx1oe
PRKh9rdtfUHnEyhpMJOgMj9xlm0n6D2/nShb219h9dsybAYAyjcPc0vSpNwE5h2dFWzkfFqgHWvA
KxF65V9twBAsguBrFIcjC6+QVr2QBAs13LK5dF6cdvfIcM+/DPRzQZbFiZWJZ5a3/gQriiMyue06
s0YJAcmgLudCgz6jvoxOyCNywhWPArjnEaXqJCD+7dIDG47l3II4NwHwWzlDCyCoQl3BCFUL2cqq
CH4zhdtlkUXgip27iNkIUT+UYVirFv1yGvY3JjTTqbFshdgQi0rkMGSuB/rpppJb05Ax2VKm/soD
p4CwS7FMbnhu2DbnoHs0TnZcO33mqXSnsxSxlCF6KpLPRazcEQtC/+92Q2zJQEgdnRT4cGht3ozF
jWFPJ+hJ892YYLfH6HjT9eGWoISbEeeKEfa1uo1xdvqdtR0sU+8k+5NDnSAD7ahh9BNe7e8iBJ80
pe1ktAHwBdkaTiTl2FdHfTA31ljbicmGVnn9hmxAzFYuthWqtHIQGAV8IPtevvUU+nM5G40zPLXq
rLTXLFXkBTzmS99gC6C0np3SHsaxyEivId0Fx27ZdNs3NZHTNAQHNxtTHqLwOM9u4Zcqd2yVuouH
mtb/zBL0AQikvNxLHUxC0RIOUtxD8T+aevYcEabJISJZ2S1FwhA9ok0Hg3kpBfrMQXSJEDAlRENl
MsWGf3fovtJ1SKM3nNtmeOLyZin8+6rRugKtd/bwGj9iMiGexGOslRxkfvpNXN2D7cmInAKZ5W7z
m9jk6jukcROR5ql8cJviHVImsTvCWVMuYoGvL28mwN5to1VacpofEitviTe+NwXUMvZi74FS/vB3
IFKUmHDLEIJS2sP03owQD5qoT5pp0vF2W6r1RE3xH/Ctq0Dzr9FKwA0lM8o+abjI4ZMlByFrK+vk
UpR+qHyWatTUHRFslaeLos1qaG1qLyKlnspDf2FrfZxHz43q1Af5/X8Chh8AINPGeuQJ/ovuczr7
HwNX+Yw5NuRTtnQu//FRcodjNze4RbNm5tH2iatCx2eiE6pvOt9NqHFMivKxzR+KFQPA2ni5Sxsk
fYIiayB64gut0TbyXXxs4ZWEECrl/573JeIuG16ZLgN8Xirmibo3aCuBKZK2dircSlspH/OzcEBk
Q0WBaei6sHQjGcTpnV5T5EkPGGCU+7VjduzdnRYGxbITJYlQHYRlFYDRFCBrQh1/u2bZmosCj+Ow
ji27ehADfJKl/Oe2tyTadMIHWoRwRpkEjDElqgXYQc5fIN4rioVGmpPMWnPF+C3tZTRZXuFJqxM/
1/3b0muQAY8yTkqXYsG01sAJgS5PlLZcaIP+b6TuWMVDYyip8sSM+qAJ+LvSQWWnwlk81L+wrVVC
M60/dD2JMq5QBc9ReEid/k4EOQLPQNgEwalbA8LBUh0UeMDxDhIrO36/rtf+7FiG5RxqxxMUsw6f
MkzTtyzaHD14uq0K4vCdCVGaUbaAeV5v0ZavEY58iMp/qBvWaPHF8xr2smiptEuQQrw1Y8t9bw3Y
g1Wz9vIVvXuaQaf60csW4zEcA3Wr3ljC/kUiarcBd/5G3jh0aQLsk4hAXieeN74nhVaMpwpCS9wL
MzQ1kvxVEa+JFWztiYKAP5gaU/tVGvizzuLGT+NzqGQ/v5deflMy0LOgdFdMKZOMpzyrCFY4Z+Qz
deX2yPfjELQdJrX4Bw5fV4nj9HovbXLbcnixkwtrK2drcjEtcIf6Sm+MybFE4SV28hUtjyyoFh93
A1QcsNxOJmHMnTMv56gM2JYLw9HDenop5KCO58AxME5lX0hVD6M9QXER9lXfIlLRziQMAApREyzo
xnjBJUxi6q5YOep+fyPhjkeb4KwRmC0syIahIy6jXLf+WospIPWwD73NzUDh5zusjYG86LCugvmQ
cqmd9yu8+Z7n1e0RIewaE/+wu9sfpCit7vCd40rPQIjP8jayWbhJ89cdQV/bjQ/E1eK4CWZ6OTie
jpfEPw0gzwaPcq+ujNuW60czoYoCafJu4q04J4c6XHwLp390pURWvO+f+rGancI4CRI4cYydT9A1
JC1mFAncrHpCn8htYxFQlWv5rjuQfirhsf8hGYk7SfQoFtdDGh284gUppLE6ISWm9rk7l3P8khZs
IWIM6bSUPHF8+W8V1saSuH/Jv/g7Bd5G/1Qu0Wrrl/PbJj+WmRFB9FuCkFnjhnljNa+Zn5IN+NWP
KiEt3p60oD953aVbEefGYCgq3PKrJJ/XHeUIHQyRB8nGqaNN5k6G5/L068cKYMDm/6Y7kebytnV7
j1WWFDm172BFjzGR/V9SuY6HEH0NX/EKi7Md9gRfNuOUJTNpnqlzQQpTbI4RIvSCE6XswXfkxo7e
UP+ssmVr1cJYU3vcl6gX41W0HkVrJ9h/2/ZUIydFSXoDblYvV5wO+l6RTBQoCZLEHEupN0hKg+bi
Aj4Zp+Tc1+GgOT/GtQY0aINz/JVlehNMzQ3nxqEGssu5aj9+K9Ta60pihIXwcvAzpYdcGiVTPp5O
B2rV2QUHpJZ/v9fvAp7f0lmaEwlRoEfJE92OufeYiW9VBooLRcTiE87+pqIXMazvPY4GIZvcA/qa
2f0Q7Vzqw1mOGeCCMVQwEPH8K/1rW+LhbJ2+8Wv60mmG9eZeJzdejfwhw1L2yCQioZ3j2l/VExSY
zFQgQnnKGLeYvmI2OpAkDbbGHZzh/iFUZntXjeGycKlpmL2+ZNBBOqESJv0I8pakzUKF05Fo1pGX
vlsnZMET24EafAY0dAwuAuwc0HzsaoAgq55D2KdIIbuGDpdisOoDcuvSsXyjxs3Dp6x3vV3J8KX/
enxcpFgecRZ+wkKm3t0IBVpGIumptY3Ct+QyYfrZnGjq+Jka3oGMsdOvOSz5kE0GVKI+w87KBjqm
RBZoobNu2hk7RRuzNucwjdogrXYxp4H4ptO8syp0VZm7bkaKXu27CvglHa+IiAkzkY4dipHNjAMa
mOfeHYRylFdv89fupnTlAm2zFGbfZpeeXqNbf3yYuL0YGWVnNfa1Wf2NSC8zPjt+xzdocbOO6Mn+
K/LhlFYlyeuvMVQGCsVio4UsG/aK7NfroivCjdDb4GWFaYPTPxrcL9jM7/D3MMHXatfgH3dwJztt
gdCni4Hizi6bOnOme74WYwhP1BkDZMtFw4VMfhi2KM+543aYqfsvQTLTOCvCO6tSOMBmh8D6IZ5c
JBpIWTWaSbE7+fGaYPS4lYHpGR30bIilWcv6jls6R/JrTshdHUyRcnHaUicgzayx5QVpftqptjSb
XmLB7T6IOY0Inczi/72ZDatd5LxG0B/E59k2NhTe4yxNGdlJhTimDRIfmya5axcRdNDqRPpk+6sX
MWXQS+ujeIsQUgLHFxvMaa/bigZIXLpfseymFpy2zzeUfwupzXmxdDkpEZrG1ZY+aze2NBcSqJN/
UXA5r3CkRYcLGJF0X4L+XRu3gm38zFaNrRdr5kQSvF6X0qh6JkNm7sRRH4O+LVK1Db3klCLpHsxu
uWq34A4u7/UIwFuveMqc5WAhVkqhSz5C+7Ly0E8kx21ofBy46uWVkUvh9LqUPMj2yvAN9IHhdaUk
ss81L/b2Oz7y6avpO9NXiNE+SVkmOgiq5RHqChdzreW6pNznO9inyB5v55Abh3LvGvAn41F70woR
0Up4JjJZ+xrYOEA6+8Iortm5DCEVQ/XiVH3chGIqjGG/sdoScqFUrcN0Sdwv8p5ymvKJ9Mszl+8T
e7yunPTz+Lx90JAFFi4ZyP6qzcjUsjd8iWS1AAtpDHyOrwKCLl0542FsaJ7RaxAw3GW6BkJD0IzW
rSxXZv7uUpRaaIi8yvzPjCc2iwSAkcMJwIrzN8+4/xVgzSFHo3K+KLBnvGLGLl3vRgKc7VlAmOIY
L4w6WWcE/H8SE2DDXjYSJUYyIFX9LmWp6L/+A457/yKe2a2/jNb7LeEV4ngJXEZ3zAhzjBGhQzCp
goRcent9uNcn9gFuhIAsrmra+dtCckiON3DWSaqN5+Z5YrO1EJJP8OVjIaE1E872cG+dQl+KeCCw
pjKvh2rXP+XE6JOlE7S+B81WPNC2dk3xKsMk3onsqlN64cyVZv24Jo+3TdD7Y67MydIxC9sLLb4L
GtKrOASZd9OT3K/GjynUDzS46XH99CxTgt2l661f9gW69yAmQUt/la6iGWFi1FBnmfEItNzaUDv7
sIfvM0Aawfh7j2FvRgYgBzq30XSBuo3TEyDH8OKSv3HFpZOHvCpuRy7XGfwpREKT2idYNJ4Bzrg7
AvGybY8FD4GyrXraxklzV/zJTD3BkiQk8HF8c7QafdlPO+qL5rCH+3aE3kZOTmUYWLGrUXj2h7/L
kq+Lzt0ITPw9gFVUc42t32wiShCb/Gl2ysheYOFLcHYKYFiwexvk7lGvkVkPDxmmKXgmqtBaLs3/
O8jXDl80YtfIxI/VsmbIKr7tPIocvddYNtFFDyz2QEOFq+9ihNh8clR1jMz/MWrzy8VhswFxy4eH
Vl7Ae4/OwFmMJajujSg0u7S0khtbD9PLo21ix4v5zv6lRZ+5ZFsP+y3Jap6dmD13r2ZT64S8VeLo
et4shM7JH1WrcvQKigE0MhGGDdqDzfQjQmcOvpxww5qAgvFzcQsf6ZPEeaJfntFKcsf/ONbDWzQc
I801Am3QESNJyR54Xp+ZJ8mO+mccnCswg0ve+DF8/lRxVyRpyS/qGmTv/3o4EiXcaP5Ev1+x2iGZ
iuHoZZ+A7T4URkRG60vgj/1dZN14WJcbpliFKTBH5zoicB3kNWODtuL6dBcNYTAZ7JZoTAlqPsa2
7zZW08HXwmZdtw2MyM8AblFA6VlJPFvQudfoYD5sENgiL7BJyajcyxbUz/BWKdh0vEB2Yx5An/w1
WjXtjZ5hRc3HNdIHwPcADqSdE1cxWf+KCHgpktHMS1kCYOV58XDBLJKWdwL3K9eYmmx1W3fZtraR
rCJo0sBgxqTSeNg4KeoVS1e1N+r46ASyVf+MwOlVAxDz/CtV8COzJXr6tnClwt5AJb2izYKrpL+C
D5m/ZGTb6bTHoXl12QKU8/S5jzkyCl22GgDJ1XAjVwiD8n4ejFiGcgsdw54xHAsrSJMgFOwM/M4u
j6qjzRLELZVOzeeBrPVwqxhqbYfSjCMILASjxO6br13PiTYz3xtNZJluOTdZ1iymEA1knl9YtL7B
CDTfMT+/HGhL4Yx5FSggi8FKYVOjHBAKWso7RhrZtsy2q8YloTU5ahXT5hQlIDZoqJePez1FU2OQ
whyqjlNY37CA3OxsAmMjbWs67TYXofXCGyFzUSBJhiX6+1Dv3VxnnvejW8G8AWJCTCrD8axgADbV
bdvicSgepa/lzBRuj9+uCUUDABvnhqCCELFqTGfmN2KpmZUPiNss2m1hnMMKWI/girg13Y2XnaWM
502UNC22GmEzs6QoY4LrVvSAURfcaMM/y9oAcPbNdtwnmYhpvCjj9gZZPCSC058qcEYTQ/HwRHxE
J+Cjuv44cxxV0F0rFNVRUxvTEogyFBl0zlop/nP4d7FSZkQUKTNWWKnvD8rRtChw5KSOlN1JBcFm
cg2h4D1MBr8jJnKuGigcY5SVUpA5nwLCf8pF1tOmDQ94HCfAQZtTr4lve+H2aatrroDGl4Byfphp
uCbt8s8y9VdXkWSb+DvWtcG2t5dxMbrkGG0N8aO7tv04OCKo+798aBzTzcLdSHC+JzpaviuVhjBF
EgP/E42ZHB6UOvW4JIDrdh9VaZYhZ9AIJCCqAxcZ5aJV97od1ELxRyr4C2BZg+t1JoAjMuxSv11M
QZoO8Nc8SuEo0pmfWBnOYemGKazuXi4uWgvwhmfIszw1TKz9I8UWY4yGZH6C0yRpcGKnn2Bl3GtE
blm0vCyDZ8OLcuJGY8OgFDvyFh3lpPagxlx1u2/+NcFblcjU79L11/mNHU/9KYztGfponSXOTeoq
mRw0KHtPsfDL8RnRTP7ZQ9oJIoHerx7/m2AUcvea1YDFcCVFdYubH7RUVmnHSvoSWALycjG/7H4M
vVkvdIWX0GcQLSO/m/wTF0wlEnMEp0KE0yr2O6VVHidQqWo6uTe7jSAl6gOsMn0M7lPcsBw376xG
ys6gKfRL3AExx4NaQudNY/TxPrE+Pw8Onj0n2DI1j7mBqDPbRE6g3XYGjAqT7mHtiVtMkXLtO8zK
X5e9XdLx/7PZTOvUZBwkcLq3IJIpMWvcjhjQaxSRDDTkWpXghPf+ZkcIQTPyTKZFo7fAUDWfU9TD
6/brmsYAEXci40b1ZNMBmLFVyGfZrSCDR4KgTWKu48lxYL9y2/fkrnBz/Nbf1krScGAe7aTBK+yv
ZUbG8dRKUFL60sPQuhcrIDzdIRG9qTeytpaBV/OUWrHxVnkE/v5/zmr4FDdC9uhx3ZD71ehi7rAU
FOO/4F9Ue9KUqOZvJlHOdZ4oUtSwDgcp3vF37U9EDzYI9PCDYEqdgrmWTLB2FX01z7SrGQwY10Rh
yzOkDYFaoyBwReBTyIUea5kRxw2+Pbda0xCT9zrxYG8+xnf3w9NeyS0vthMDH0UGOCklRvln0MbA
r1PF63mwtsA10sUrpkUv18epj/zsKckX4ta9qiklV6fkwFioCu/avsn/QxTB9i0SLiDKL0zC0oE1
2cCYVKh7yTRm19RPwzgxC6N30TRPBkR7VCm2264A8KfM8T4HRfj+EiOVmDaoDDSUy+TzB236zd+I
QTKBksrjQU/TUAh7aIo8Od99M3qvQZ0ffv165awi4l5x2tirsdgXltFP/SlSnGW+Ucs+oGO+XeI0
EN+chjvqn0YMOJ4MQzGH4zcbhfu3nNII45Z0Rfih5jCrwAuV/KMCflcpl7FE7Fyavf/ADHMfLali
9TYavBzdp5ZE4hv73dkQlkdHH5E54vilePtlkpOLhel3yP7wV0EmJABghAe9DdBzO1ssHEquT2Yt
MscwDP+45psqfcM5mfhvRPZ1OXgUzaoKl9PQ6DX1s2bCurrfoGZqLIhf6rRUfdRTiLlcyowP5QMv
sEBLZbUZr0MhamZP6sINdZU595vEEqthTzWApJATUxtEd2zF9KlSgGhS/vaVVpbVIsGCcfXbPirU
3Y9YR4e+5TuLO/i0bQvcEIeGsZrXuvhztc4Rcw26OSbXd5trVhrOP/ZcsCoqQNcBRsC3wSI7RUHg
AAEfFoCAGYqIkAfXqW0ErxO3e9PO0eMTzlYwu4vm3hkNhLPibeDKwdp6SyNWSvOrGEMuPZbOH+sF
a4r+3hJzNntGjERcf9MfvTMk+K3BNnmedtVQ1u5+ULB/cmq73aF9s+x+pIFCFhkYQbDS/vdXRC98
WoIlyZp2T9D5ZND8FCsdRvGyeeP+H7eUfCQth7/ecPwyiE1cy6rv+CyX5jQqFiYtOn8ea/N5OwO+
l2xOIfdpo3f8eV/5qWhdKLkhXkc069sdVefj1vLg1PklY2x/kJqTs+a/khhtKdLqiwZsB+RnYu5h
fIwPXBlPmavO2+ujgSkCsbQ5Gj00AwgbRuUVpOl1442qjjiDp1Obw0uK48qRJWxbhkWE0WU0jlVL
XvWonAOSucvHARpVRBu2lvPToIBfJELzuPNvIfq9EVk5rX6J65rQyu9ITbsjJuvWFpTmbBcMLxtm
CzzyexzbqIWaK+bqKCdqntugc1qarYNRlvb5LqfddA1nEbLBLoKcAOHmArSgUlSQpC3STp27EPd6
RRDoUxVfFNMCJWXu04VRMC62d3KOrwVldIQSb9dt/0YJo4P0fMzXbhC5nrAo8DgxDZL0tgy9pMjs
+SpUkVLBNmgHXcTrabwXnhWiAmHlHeiaxZasnaJlb0kD4O3GMcDjsRe4dDGx7gsYG9+/qDHf3mDs
t0B3+dPib845a+hSjtPSMkuVkujxaY0A2BtYbAJ90+35sV1Cmc59hVwqJP6fVAsWz05ifWnAQGg2
XoECjxRcPjJbwf/DNwjz6Qh5lm0bw9isofkCQVJiDmkEmMewlFVLVAu89Z4RLsOuA8GvomVrRD3I
x53VUmWNohuV+W5MjlRWXxS6BClRXO5DIo4jz/rsAsPryLKrJDVt75tADVKzCW9cHUOWF07dLdrZ
eC6vNcIJpjQmv1kYPubpJ9rTNqaRb4T0vGnDVDxdqFmuUK9WAP+8wVunniKwPfv+DSiKosP2ocwL
8KLFRMPDLfu/VfncmT5Orqv0q/sl94MSvvo/ZSFB2ZAB8qJRZZbFqE6IgejntcYnBjUPE20gw+2D
xFIqWHPFf0sjPo3fpBjbtcEJptkhiVT5Y+8j+zyh7nVfIi8WncwJNRYEPj0jhZfoVDxqEU5/KliR
OZdgf18DKDXjN3Wqxx/IuB2WRXHnAaDgAyQP0ByVXlMarV9/1c+u42mltO9uyufL1v0wDRWwjunc
T5lL3eFNMZiwyMnFWte/gWKTI6QiHedBMVw5G5tkF741mIWdSX/gamyAXHIg5pvicCI9tPHDRzW0
DtuRcKoiOrkqSTwTlsWzjZGPKSUn0zfAj/a2RxrWICnCykj9qtiYfznXNpP8L9WSoa/1StRwO886
RHKwdSIx1G/Zz9cmTYin8/m+MDrtNjhZSZ1ek+M6gYCKjVGdZzBLiMBx/nVwukkZB4v0iAa9yxOl
jnmXgClTZwtsNsxW0IKP8rnant/5dXt9tCiqwwqUIgyzdCbqXwGJxF20uDmJYG1X8CvADZiBf0kv
iM/N15QoIzxUWapH5Qlr9MpfvX9pYgRwoYHHtF/f5UsDULn5D7Fxv1m3J0qXJFh31mBQsPtMOm+3
1x3nsWD4H23vxdd8OlIBKLGprhQEFz856rdQX0ZtxTarbLmEp0j3vUFTAzAeO+cj0bSEj61dBA5z
jZn7ZSi64RvLPPDrFF9DYSK+6jEaFdT9/jwpzUerIad0JtzeOgsoxwdp9VEfN2q83UxEHfjEMOGN
TJOMvdyxj05OSwOiB1+Ligi8DcyMXS9d3uDmTF+17jL5Rd++XtD12JrzLXnJRs5MtX15kCISZFDp
TjPIuQ8pz+a7piLmfHyIcRAUCZ+TCJtn77jsMuxkC3i/Lta1PawzG3Km/7zhIbG1rd3a3/B7Vu+X
X73B4I8xGO3Bo+aAc2gwVKX8C2RfDKea1AraOLXUDiKy29nthkz2aRjapb8e0j7JzL8jnQiop3wu
V2I2MApPgLAtKnaFgH0f70bbm5HImPM4G9Vn0Z3FYYRwVfIuxWTt7W49k/j/736R9aRfMc6WG4a3
IhP/lN2afvP64Sojne0+eQKlK2bM9AIIhde751hCrNL0NssLdUJUPNWOCdJ4KtovnkhgvuXw40eS
GBl2uvJijzoL3CMRN314tLvmk8JW3okbf32T6v6iwt651U3b9FlmAiVthtbd9Av9lhrzrEIUIrTC
TjzxdttIlsCmR8FYhK/vX/nMYvi0pYqOGgK5Qo1ookMnMGJUEkFlaGl8wCZSzxK8SS6aEuN1xe9n
AylhxcHh5FFwdAB/4IceMVR01VMMG6yjT9L305PR6sYYrMi0sHVIgDfVYXPrREjYrFEEWeWFhR1B
QtHbKNadLhN5sYi4/zUzmmfJs1uX1Rea2EP/3ojJhz4QfHe01qSai9xLvHX/Afuvr434w1eygr+z
GpctG6IRr97uk/0yyES/9RAKVDoCuu7P9RDyKQcAmzhFi44Nj0e8zE3Mb02v8uEVXvfF4RAJQzji
MUcmRVia7/d0EbTQGCs7jiuEuzjRrQVQMQDYGGpxbOhy4lbm0nnprWj0xn9mOCxLPuDcRVOdCiDQ
mUm3ATvYYoOdV11RTP5KhLLdVS9Hla/+75VRUvMb7z9W7YiPkPcJCSvR/RLqZINcQTbIVRGR5lEO
1lU0JuAacz+qwyQE5vafZw151pU/zU/aid7TkPZvdfx7rvOwoIOKmlKKlWlow73PRFIJEzuOp6SF
BUlVvmXfTDI0uLFlXxVewHsR1o37jx9hNdCjEhmApvC25aFYousCFr9GsFW45r0CnUzUtLD6d0Vy
bJ5M3o7YgdSoCGGEyU4UOKX7yRgp+lyAi2GTMz+ACUH5ysSu+xtzR0XZ90sZtSFZQC9gVrU6FJoK
F7d4UkIRTbTeF+sAwszdZPHoUnBWPlSU1KUdjsBXgUjhd2W/3lGix8hdPQtzRux9nNLwdus7DdBA
YOnAhTaJlukaNomGeaWuEjVb9e3X3BFjCpn7hSEi60UQOVEzHaSLexo2oKHEf0kQ+M00Mo2usdEu
ZkgKuJFbT8pWPoMf3wmqntjX39FQujss84F3FnFOWFwuSgkMH/sTx28kGFikpSwDeDcg66MWKPHr
Whr8h0shSFYpqKwA+idpIQHt+j74xxybicZWaFG5nUo+pwA9GmUIk37WyeaDELZyFsP6jcAZXvKQ
ni33J39OqRxB9Crcr3x6XgBt90jghaJ9GlkVli0fmMYvRxZ15SfYEoGQ/Enhn/f50KKNuDRRmSSd
NubnyyTa8CitqPLGSqdMcys4NbqyW6OBx0SvwSaoikL2ESN3LLeTzn8HCMKdJeeZPXLyJj13z1uN
8QAIsTx01yhmUZIhkWrITRiD3TLaoquTJNKMF9dsXmkiuayWLV30b7ZA3OAo6N4G6HyefcQqZgPO
lmnn6xzBvaQOwGigfegP+Ns+MO+HBiLwE945ov/H7zsjAQ5v0MnHQfjrF8SFtiGtofbssLdeI2W6
2Q3FkNk7DsJ6IUFZyilP0FU5P5xE6jJas4gRdiPetXtIIuFPWsTn0yXqplAIU3mN7oGdkF0S3Yl8
VNqkA8UnEzdYcyJf2yIIcm/eSSOVZp1GP5+dUEvdpcOEUppWUotrW0WETP+Wkw9648JbQk3jrg91
UIK8G60gOJaqEoMr35+Y88q9GIdcRfyIHgnaYT48Kg5RiFHRMTEThbnonsfnZlzTMHqCcrHT8B8D
JugANKdWiZg2WvzKu3HK0lCER2o8OWLIXiFRARrH45z015U9ph4ldKehUX3zm10BV7PrqybT7Dbn
pgQXZsC9SVW9cXbbmkTD10UUA91LriIXtqRehzrpI91lOazLassWLH18qNIcxliRPS/WNRixFhCX
dSbJ+IbMPiX48SscXM+B1X9llvuLnMc8jxkN/cwcwiFnVPDDXkAGTQiTAb509q+FmfHGGB5fMKLz
WGCAQ6jCkAcZ6LBtWann+gIt7pK8RiQu999IOE1bAapfkBaR8Km57tNofUQJNZMGFkjBxgRPuXm4
Je27KN+OwkRBj1y8ACxGrah7noFyBsbMQ5diufhMOooIv48EA3sxL9HDTNLJDOseNDKtu4EbtAUy
1hheF5DBjqdaKNMx+3J1HKmXmZPAAi0tIFLYylwTBYoAKECpAg6GCf4Wy6fJxz/m7MEspNox+Y0x
s/gngtSUIG8pUIXYvbowKVyqQE741+bLtWGWm7GCSNx0zzoLwhwTg4K7doO0LlkUAPMvBFU0UUAt
qf4XTnyOJlki0z5WgnwDF317h5zBKqZI1yv0JIjdCGzUYgSvB0mpQcgttruuiA1lVATYXmncwu6L
dVdBjdfPIQ0qvVk35mkQHBUtvk51mTC1/A8VroTIi2G0o0YZ5kU0TdKoSOlidD/0CPv3KbSxfdjV
Zb05F7fZCtwg8uCp41Z8K5J/olkjh2wffe2z4t3jJgYOwS0KVtwcEtk5h3sp/lAmaqxlbSiFZ9TG
dIF6dhoAOTmtQQM87zE7pS7OhPeOBemlhYZpCujiL6xjk0LTx7k/E+syHtchBESvqLwUKRr3EhLZ
SGynpgr4QBlAqRUkH1d3tmZ9I5bLSLCceAfOpbGo1lSx/PWza6CTNFDmQQfK8xb5URAnb1pUfTfq
ialDe8qtUqbIVUEQjHqd+wDGCUfxlBH07nLVjbYlPrnGD0S54vExhenV4vdNcEe8o/VE5k572cc7
sDIAZlOPUGW6uRxu8WzIMin/vT7KeQYmdfaSewpKc3ITbxd+4r1CSu4imI8Jz0X5OXMYZey2Z0+S
NSJHzSfsldQz+8H0TRjazU3bMXhkYzw89Jize39VXDWiBO4/BG0mzxTN2N7Gth56YA1I9DCgNX9x
IsXSahBVamZoKwCiljsL/u/8V/X1XHgZimi23eLoRlNlHO7nLd/s3xTaAR43dOElfMjX6oXf2RmC
aVBa4+9E2QT/vQsUx1nByaq9lgyr8GZt10P3H9Bztq76hR5MXrn0itb5hxDWMmys+InYoWad+vGV
yB/ox9+tpgj6eqWCk56KACcvDDs2S6UKyRQ1LKkKMXViRdulesR51L1/O+cgmBtNIrS/rIbg1nWe
oCqcqHkb+FxwDdLpa6HD0PjysVj3qUSl6dVjonwm7OWU07bNmXtm1pn5lYD9z6nSwsSuy7Oz9IMG
lm+n0xBAfOSZUxRWVTnwjLM59kqGWr0S5VwA68/RBgy91V+XgJ5LoTpe6e8J6fg0WaFhoFjO19IK
iDvNP44WOsRB8+/aVg3d0krWYT0H0vgZS1iNK8xMJZx+DDZFmm6F2Eyt/cRJZancASX5zutypO0r
e2aGLvEW9N2R+2YDC46lcM8EyAqJrdgwcwGjfL3nTzlQ52r56t124QjbVMmaBatcoL6xkCHVDnLQ
6bWRXrEudhBwmk1IJO7dQQgPkD7bo1HxPJpxXRx8hj/oLtYlbY4FXszaFdvgnvMWoUJcQh92Fw2i
LqZvmYfm861S9eSUwcPcEoWVCaJY3SLDwYDUIgoys4lcEl74oc1y+uwB9t884WXCo9mgjoOfYcr3
vPOgl2wNDggaMhKFPPZ5F7uRhvDNI5miCa/utvjOUn7K37dLnb/DjRE3W0zNXIR8TUCBBuUtCbL5
MuA5yqJw2RKHRHv8u7gjcHmGg8PFgLmSii8RJvt659UdQ4stiRlq6r/FwFz3ALb8Qz2hRUXuaIwl
KK3NWrlGqQR89yAtjGGTpnkjRz+mvrvO2sRYIv8X/WWQwu8sHwkKwkKUnN6/xYUbDrmRx3uAMGZ+
a10tCKFCWpRYI+sws9TIJusWT+aMficPZNWwGCVNcvIbiFKQe41DCdVanh7DkwG7PHoVP/17bGWo
MusEcK0bOkJBX6/lw81jRqMrYTT9irV9JT4aldWIveAveyYHQQNjvT49Rt0sZstYlYkWvFXEBK++
pDZOPst/gDpDuLFB+WRYuqZfA07xm/HsBhystYg9Se4JJg9iuOtaZixAQ0rdX0e0bNgya4tMzXp+
8MJiKI8xdLBuo9gBL6bkaIzKYJXK/GSbMXIkwH3Qk29aOmhanYDSBsbpioeoupVR5qIMj0n6OrFW
lDu+ZUAxCnj65jCd5PK/4IGSkyOQRsunCYGUOxWEE0hRWs4M9g9AzDnItoxJkA/WNL1i1ZR3fDxT
TtifdFJUG3kQgu69Koqr/Tg4ZtMafjdiYWFaE++i+8l5mpZK6imNXKm2PVcRRHGoeszeCFf46SvQ
jK9oqYu9SGlSuoVzm7KO+LuLlXbSQXNplkmp7F6cr6ziJ1zGr+7PP4wvrvt5j4ZiKAlKbA53lZ7h
USZ1hVF63CPxUtawtCeOtgiqnYN+p31AJDAWAYIXgWeR50l8zfAV/XcnUS3M5sMWPrlA3PTO+aJa
H94Y1Hi20a4WNIPEcJITPqp1gKWtdggB0/VXTnFkTjVI0g5WfuX8JQeZMeRpZgZZECW4SYf+9bsD
59AX2UhCMGDb1yLpgsHGSYvUuH5ymRtnu9cOn0g+EFeKdHcnEd+I7YXtvQycCnWx6aEfwlPlOa2X
LGM6GsXX4qDaH5Ig9krxqsQpAkLzpGDjpThMFT22TK4Wlv8uW+dP93Fu9CS4u3ZEGpwxq4ApwYbf
zKTFc/2JFzRTTqMf0CxcUsPCPFG9n2N8+hvjGKnIV5mtzZkXC0XoU6oFTNE3N0sQMLV9h3nfJK1l
BxBxkXS1IeUNsbA19PkRacyfOorimv/ho8ck/U8/MB97mCa1mRLkKut0RZ9LxbCX9xf/Kl5+spjm
siIORaoF3LDZbzph1vh40LONAL5vmPfYC4qp03X1rOK4JlNkD6/O7uTtg5x5KHZ/rwsg0kQEVI5A
jg7dPAIEzvWNY2H5keLNf+szGEMpRQHHmZu+OEmUoMvnPOu/tXzEHH01R87WZy/YZB9YnQbKpl2L
uGa41kXpg7YDfHXQu9bCAqE0i2tScTo6opB02tB7ger4Z+V5m3e0MOy1RNHduY/2AsED7kdsGt/n
B82YryKAAcf53jwUDuUICyZnIug4fkSkzT6IsxQFOj3lpBJB8L4nf3dSu3xsfT2Kv+YtOiizwy/8
XGI5Wp+pyt8BKZz/hxhQBzhNmSenBQMPsD5flsF027XAimhqNUt1u7X4MFkrcXgQ6Q07zAG4n2Oz
GxeSaQ5fILFlx0Q0rOzkwcdy6yJwUOCDmeWLWpD2YnZjEEnBpkYviUZSXqTSyxQ1hKWSKyJbXBWa
ltjtrzBwAQic2OHJMm7K8cjpy/LQhoVBgB0n4tB4z90PkBildHRqJCSrI6Gmkw8E1atp/Z6j3+4o
Zi5iCyOf5qFn8uLi2bvK5BXSXtvvNSDvpCs92qdmfXhmwfmXTfuh2DEhUwoG2B4J9ZnjuXpCGaFK
XOEeQQCnocHyOvgXfo+XuSQ5gnGFxeYMgJVZ0Br2KT+8LKONBPnmnC7Us6pI4oJnX/uGJw8uyURZ
pMm7Ue6tb9JRTsoXOIxbRPSmw4EPSqvNpOVC9fJGZ1A4DHwAIGZbwbZmqnBPM2y9RzqUjpmfo43r
Rnl6DMcRxBAJy6VuJkWkgSUNtPAN4v/MKNSmZLyEHh5PH90P9GYMh1BuvIKK9Xf6xm2yzp7O71Gj
29SKxn0TTvuzLPKV5/33vcYAcHSL1EatlsOx/xow4aKRQ9ufHoAFg155ILdapMfpsodsHQavR4QV
jCKzplW7p8pWADG3aBw4e31dTfRrFMx0ABpKnLL7aseeSEEPD6mdcraad8MGAJi2qz6B9oMkmhxr
uotGra3G8lyUKIZ/5+E6gmvUoPfQ0vZNuZEMAKODEAqWrTY+hiK2ASHJBmFdZ1kye9io3DC92WkB
n0gRHuEmgTf5wClwQTdIXM4osoVl5TifgFDSHEfAZqq6dIrVZM36jdjZKA/qBQxzRRNbP6frAtY4
zcHZs663jOOys3DkP7wrVghvF6djI+Y7gQt4CcfXzbRQXbevEBG7VlxJdsAsi7ZWXOQ6WWcBPacx
8j0IUNUYfurg1yb3V6KsGUfljb9THU1WmOLk2vMk9ChEvMZ4rykzL6QG/B4FgkrGW2/X42MzGLG3
vVG6Ayj66Ohk4/TguMGQH0DRw1mLo1GfcDnOFkAdZI3BoqfalRelx1kWcy806zBYr5v2pc7j9kMF
lo04ov9zTw26u5XHOIXkAUtMoapW9odiLOS+dqECceVqPv6ZBMFe9CCZT535BjtmMHVmqc2PnlfH
JQbUxhdvrqiIGG8dEWh2WnBiDLfUgsi9C3ShhbFHdfaFV5Vz1JZPUxgp2ixqaMdslwYNNKyneRXq
EfIUpjsl0rV/U9L7BXD4Qloz2Q2LpBcUR4b0pYys5KBkn80b8IhNVBi8F1QrkzzSZh5ApkBguoAZ
ACqT7rES3MTnkZ7ibeiEAiVxEaxil+lsMpYSiI+hCpGkqo7COCZdv7Mpdj82cBScZZ7cz7KUISvS
zu5beJfGHAHdePndIdPVKHb7pS16wn5FaSBW+4Gz1rCQA6C3xBpDSIu12tB7sYE9iY2l9ecYWEM0
uR5TDQoFuaD+IjU1zlXTdhtTqAc7WmGnxkREI0UKo2RnNIBUNMzwASLrme2iF9sYSeQDqvoV/ujh
vEH4qnnnM4KW/IFVl1AJ+B+NQBJVtA92du7fK7ILwQq9yMWZ8uG4pr36KsqrK01c6sVaXaCrqBJm
vF+1DXJR9SkpV6k9M6e26Eu1fkmhd5yzUQEgAHEdc8emZDF+zckW/F74y9XtSBHKSw25rVvKZ4k4
vjeUqEK6AtYL6Do/byx/EbjP4EtKqLgZ2iEk5dKa99kheuiEgyGwEq69GTdtef5jbHQEfd1cve4I
G1IILbWxiqImwbrDD7XJoHK+c4P9ulJOiLh2VWQDsYtuPqa5gTsPShb8F3yCXY6XIhrBn1itlOQD
+SGv0nD/9N+GxFjk+S+xTogsqUxHB+G/hBCj0mSgsnBgFmg8MGPiHDr0yhTc5KbXLEAPPfb+X7vB
rk39XGFRa20jSc7mmD8pMYCCHSnx4VbwnLewGzjX2StdkPXZzqPDnsYMPk8g/m59xCPSlL6gXDCC
AZE4dxx0ojEHrSLSHDvd2XNavvlrysaNDs8XEv6A49Y1PEsUkJAdbfX0W+sPmNFjkvHTCWpKhp3X
DAnMPB8uxbpezVb4AtxuaPZXOdhmGiZCrL41q0wG26UsQ9gooeGnsujwa4VDQXu2aPgbb58dGvXK
l8Qxg+tLDtsRV05bTvzKgaLh27EHQhHSbOTsD/LN2acbhgVY7QDPxZpImJzVB9Rk/ddaTTklp2Y9
KtvBkDKPZQVM04E762HMo7rFrerVq02hWNDHSs0WlvEUK291tkhOxzSOOUrkSXEJEbUFvUrHP/kA
RJIO2knklIwTKPypXBmIEgA6xByv7l4T2uOK16/eKI5K1LTjiO6P8qurE7CrK5nxtm8PGlNipJ12
fvshlaTavSVQG48FcJ6lB4bVYRrnVRyebuzfv1qq7F4t4o95DGiDGoa8T54cT7SY0M5YxBC4uK8x
cJgaViheDaUONXSQyTn8hNgPQJQS+36c8Pp+BkbLYTW/oTPisv9Rqd6NcCJKW0Q/tK0EjzXEkuOl
AkS3/7sA57HW9r478Cx4vu4vf52q0XaJqsJntR+kHhFyQcDv+IBBqeXMzMmd/1bmTb3/a7RDMO+D
zHiSniGgbRUbOErkcFQsQdl+puTmEGlKmxxZBcQoq/uTRqHGraKkpivu0nurjx60ANJNe3vXe6Qo
6yBqWOLkBPFQgAUCC9Sdy8lEm+ekxQV+ajMM5Aa7vbjjtIZLeR7LomY0IEpKCEMXoklLveJHEDTA
q/zKkrkBmX6uZfbBMLD9NHddvCPa4pAiT70X1nsVu0u4YrHRcMuY9lFBH27T4FTkCe/2qrwkbZD3
ffPtfKKoOf6jBhXWXotVp44AKgASeafL+WGAHDbCppcM3VSn80sviHjwuEFVirsQ4h24T3DChKGs
fpKpEO0qhyrqMXvFRuT6sg2WnlgpfAJPCGKkHK3/ov92cn1z7ilqTXqJ/KMqNtJw41fLKAFuVfZJ
p+kBuGTDdYlTTKP35gEuuCIzpy4EW2U5XiyvYJie2cTT1Vg9YoVVh88lthI3aVAdTjAVfvak4/fH
r2G6wFBIildwaUA3MKRfX0I83OWsqR6fz0nDyr83+Rqkd/WoNYWDs88k2Iw78IU+g3XkHoQUnW5U
ZCs+CR7gpxjYO9FptETbitdTba1zlqmuAhzUM1226AzLbYOGqr6dbOVmzCczmp5/LW2QKvxcK2d/
a4XGuYCFR8unq9b+88asRNPAj/pQlkWdSIvoD4QTdp/ByamRzHmj9OWCMrEpfcBPLqYOIcRe4Zmv
mMjstwlRzI/3tewcrxSToQ19yoMdAmjRsbUPWax6ceeAFcgqFzmn5CMzlHg7HgGfGmMhheX9Gpkg
atMAa2ZIugVq5jlhVrX2Id4Z5FA2dMwh4paskeI2LyOpwZM63zJDx6adXM/+B57vP8MbLTDodxyF
Y10+YFB9Bz+SJwoJjY9Ts0XsiSaJODVWhi8pXiW9TU6Yjf+zQhvDh6ubD1wnG3UC1gI7iJP4PJkZ
4iveg3o8C1dlI9szLW8OoUYq/Up6Uv4bICN7IRRgrYCMdjEObzdb6P9+MIxOoouibfuyB8uGUSUx
HH4csBrdSdZ6fFL6h9cHTJqW4Jf07n5CJqXe3fNdz9DfFf/ypnY9jy7SpGygh4QP5RkTBIw04jEC
NLZn5wdNrgMrtmH3VA+6Y9RWRX4Zr/dz59hvqBt298l6/l6473O8yOluC6p7SgvzyVHg/+LxnSb6
8DxJdH6SyjBw8WFJqBrcgQRSSrPVAXbnc9PLN1gVSe0tML+VheT2DPyaK1Z2Kw3JkX52W7lEHVA5
dG/MM6FeQkM5Xwn9ynB3Y2f0heHyQ/QT4iNbtLCsLSsTmngMAZH7Q6Cjm3GeExnKMZ+ofPNpMWky
wQhwA4Zr4tVjvOwXDVWf9jgTvBPmbywQRj3m1rExuN1qrzXPRYTudrsK95CEfoRE5QGsj/X8Oh+3
3VBw6h6fUw3gmBgOR81tWufmIbQ1WQlQD3HeI8YpsPQ/d43AuC6t/YJILhjMsFwlExNw4tNCfDrc
zIKxHhtHc22trAEMrGKP4KNSoqi2Q6ZEYIgZZy5OtP82d4iOi6UbYLi4GJ7hKYeBncg/+4y5lvkg
l4y1nQsxE0V1/bQb7b6hTbfwPwMdxpKMpwGTc+iPr4oweVFLlWI2FQtKgfU1mqGWH49LCaaxClZt
b1SZF21jiL9yp7Ow79n6FhQdScVY08rOnlp80o1SfDbTuHJGU2W2Jirj6sy5DUPKRAJmY38fFd2L
mS16gcuIoYOxXSHazNSBJHOgJYevCegAA4efftRCsx2FdYEHu1HEymPFNpcXXcgoucyHaA4mOoc5
gDQwrIiFZhpWryGcEjGTjLiAA8w1xkUcyNb7v0WNs+5GJepOq4vLlgk5RjUvqyvBxeeEyiq9Nvy/
yyINqB++7Oq/GV77jV2y6OU5IFaNqIE36/GfKSpZftBMPd+dR+NIfHoJ10EDPHoTcb6tJ4AsagWq
3+vVIQyBA6vVR1De/Ekt9DqXA5mj/AwVacmjiWyoLiVi/JkZ3hniin8X1iQ+J2kqeGiaMiLzbJGs
nVMEgjsbpAD35T00vW2W4jiWf0vGYcCO1+euTHYZ6uOuM3UpR14CoA+5dCiVE1WA5ZMts4BRw/n6
p/+ezI1qsG0SdGpE41ZhFiwKOnj4Tur/SaphZlN35/yjqZOgSQnlAVKUvHVIHwlCN4MUow/XNEBW
x7QXF4Zj9IcXgPUJ7fK/9CZZQ86IHRxcUGs78NGipISpex1Nwis3oucA3f//b90ZpgvPawEFKi3M
klYtOrOHETUIRV9Eu6noCoSPKm6GKNmvUQLM12XY2ttAlgOQ86HSxwrNXM2lvx3dTGRh1y7FnOfL
r65ILvwyKZFrGcTUoJ835GnTFzugjJbNBPP9jaJzDfUO3ZbcmqXEkvKbaSB8UFjd/m79o4mC12Qu
MvSc63Ow9l5+V+pfnxMAnXlGsbEBM0YPaJv9tNt1R0Sm5JKeVbepYKqy0ho7JLc3+bMONB272NG2
vyDswdFMfeVvO37PAKfE3HRD67RaQxwxp4BdD996FZu+MvboUW2pD3nJDUNPBmUq1LCXYRyyGuPE
DRpKAG9eUd0NkrsDpI49l54u4wqBgkYSjUk/d5ZXluufJYmLIcBTfKPnZOCdrpk6kWRAlTh+I3b/
EbJAOek/sSwv2MYSZfikbjC3ZJj6SC4QjyqwRglwtiBboVHnNAejWAa+D7nOSWHGRD69dx25c87X
JVN3SwSa8EGpVQwklX7TgTsrfaV9ASvA48oXTR43QSl1ZNE3iAzNPfo4yLQcKJy9xVWqon5BD3ki
Cz/X3r37NGD/Y7xbheQ/jkXbxvanN2w6vt0SIIolNNxMcyBj+ToInJXPjehaeQ1rNzDqBAU9mv6A
ndBSXnV7wgqOJH8fTtjMoGQ6Q9xqEisBwArUJri/SFpI+Eq5WGd+vvRwLMrBEVl9NEfpMAk9+uiJ
/9vhe/UMS9+ggnLaCKiQkOIBavt+tVqctmLYjsPfEubXu0Z7csvQeSkBiQml+8uTgGAB/z+LU5/D
G78SqrutfuM+NHA6elq02EU0iGTtvjY1KplGbYrRDfNcYl52A1DGJP1v1TkujykkcqRCWn8oDGap
Y+XRhYGTMLJ/fY3EfWrDuapml5DAA/IO0fLpJK3fIzUd3/V6ixFJSZ4cag688NjyfKN5NYrq5xJn
LDr0t0/AIDZNDCT/z+5RLWOpJ4JhYnQu2xxaKOzpgzphUHWPW9gQ28Exjncg/xdTzXQnhcm2+rmE
d/YXk942dJ7n86cuS0HGLIIUvaDfiAy2Fm3UeFTEnXuLWXKkaqSsf3Nl9s82qbQ8ahtrRQTl5y5I
D64mRgHejAakkwuo7glz3L9KmWwnQQas3UEffzMiyYEUWA29Xw61/ybp5Uu1PkPqTUVaJGJMGkwa
DYuxX1qSNQctZZJHoL0U84I4YaindFdXsAOubIxcQeMUVc0Meqtj9P+GlKwSjpwtmcVvXkuRHqwg
ZNEgCd7Q86a4vfdTyTPXT0IZRkWZTE9mA1UMyia+ypUN40+/FDOgqRyahSGlPJSTfIx72yNl2UOg
3km0FFadBBH/BFtouwDcLH5NLqwKj4TYixB4rISlvLdEDwdeWcwaZK9tCTXrqchHfVn32g3ECydN
s67DqK664kQe64o49DOXJz2P5vBh1U5GS+APDE7VYlCWqVhiUqjFIb8wr+AI+5f1xNI9jMZG5wjY
2Itx/fm/i+hFNkdDti6IwaOJLDrPh4zs5zgZgEwSWLH4XagNDhiJWctbW+/+b98LnsW9XUMcyZIc
8AcBSTKSNddaO7QF0zwXCnmA2EguH3YAedZ9lS6dcnLqamdj/7Ghk6lHpjvYYxIPECxiV+9YRNda
antQyLu/s4vZrzWVDgbiKLLnmcBHaeRjdK4K3hrQ9TN3sezKn/2NkmnfDjbnrrjzg+E/WcTz059l
g6rS/HX1jj/G4R4VWsruUUPxWYXqKt7R5y3i2/RsYxyuTRtPj0aDImJ6f6oLtR2hr5qgLy2CjSZP
r1w694wrvsROsJszg6ZBzOr55TgZbuqPtntT4BoR08Q2n5n38J1u3DN95GaUtwacyzbl7miKSqji
KnRyAG0n3zWamZsNYtWDtRK48nlAyCQ9fFkFa3UP1cl2WEtsPSqnLCpt8la1+aEMCtNScj07P+u5
1+OVkzB298ZWxhC9iQVy8Djpd1bg+Mjwd9pp9Epfxg4J4ET/KQOKwywi9lKv39coVaeZnnFiA0r6
EXHpTaO4msQvQA6sO2wv/aDibeWA6u2Q4zge9xuwtdjtkPkEfEFOQfsXRE8nszxeksOqG9GD+xGz
cOPGl4yeFt6VtRTjzUrkoJrFaBxMwC6diMf5ii/zfW4kHSyjQUkfUa65qUzkplYRSlU1/+gBy7p7
INzcBqgWxlEK7wM0JTk3soYWW8twLnYnCtLQed2L/65UJ12qcjsNQWe+osFYfSDryzWyjX2Ufabz
nbNUKH5Rpgm/8uO1pSV53nSXplKaUC4UetyJ8wjEAYawhAFmRF3UfwGh31tJfg6VoGRGAM4kEvFO
WqfRneL+jte2VhTDhmoEKS11srvbj+h+FUfY/KT1/lMNFmUpkTKtVo8CEM2+fZrMVJdVezvWXolI
Aed3Y2lcRO+ay+39OBwJriqvK7m0gNRKEJ/qULRHgnAcCs1QCYrijqk6BOX19O5WjPb6C2SNxnTO
kGH+igwIGVHEI3GTMDFRASohs26PEmHzrFgur4cqjLSmUTzuKC4caw+uxN3TSG7c9t6vwKa79Lxq
+oA2cOovobqlnTAQBmwAMCQqKc99ZsLka8ObAFa7HBxwFrRyD5GB40xlE43RsI9aKQd1mPeioYtr
va4dJvnRiupwa4lOM8zjHB4jFW/Gu4L6/Sr9HBavf8tXKuSehXdqTugveaVCiYQ4GsbkILSepfJ6
IovDu4YAkOj5jNh5wPiSmtKL7MeiZnQGvO/uf9YAHI2crFy4hcqSIjcbmc9A6CbattqUx0KDPvfo
Jcb7id0iQDpggx/zWnR/yrp+l+YjtQgd8WEJfaobOLwQaSvqeqHnVaWByOvzDv+j7gWs+RC2AW2O
r/HmgxXDgfnoIf+YNhOVJX8ztsizwPknVLY7iQhCRFXBDAVg14nJZkvvk562KFXLhzGkIi55YQLV
b76+2LBl1DXDR5CIAxC8jICk/UDDAU8C7UduYf6n0C36/2YkpU4J1gGeq6a6CQONTe4kVXYhX/PW
/1AVnZZyqA86EtoP51RJgC51oCJ0sc2cmW2el0YtrrGpjnfLs74Dl72uIAffRxpaN4AXBPQtFG7x
i+Zzln+aURhWF+RGi0Bahg1ICbHAhi8sokEDsPRfQluSW/A8EHWZLSGpfM4KLHAQZSB23OPyhK7C
2hevUwTKtutKqi95+AgFOAPyIP2eElIVU/wx1yG9VoKqOShTDLuW1lJfEJ69R3E3Z+v72GcpGhRe
gy8y3KEBYjKA3Vh+nvYk5V0j5k6reLuNA6sde25Grz/8hrVFCTTxatQntuqpo32mWuKmxZa0w0LT
yxA3j7e+RQ77UZDe5VW2T6Njabghs+OlXvVXD3K/v9kZYdy9nzCtGUcR5fEDfm0UJDmBJOq/BGMn
vp8EEWjkdU3prVCPsCQ9CC09YIqnKkPutfO1RkvZ3ZTMZxWk0aUOcKuzv3Re63tWfj0daZK0bqyF
jYzO/PhgHkydMNWghXpoJ/sDyeqAEwBWUBif7xpm/jGege+RO6ta3XZv0v7wR+iP/ZG3ooPpkY6s
MWxCFWWkeWmfYsviAI7z1tF3X7wwVBo876qOWVvURqwZgpPxEPsCmWUzYtjA9Wzu+oWUPQjQ5oKP
L93TvlKCJfV/fdLHCNpC4+0ueqUzoP+SZm4VAGRctN/UqE/hw/X1GcB//avvxQN4Wgn0/W9HzexM
dKJDJ0U3XYUxi4BL3/JcE39Kqy5cJQg1hgkODDoATn+JQpQzdNOzwyqz2sqsZ9kXTC8ujmLHP4iT
gYg1Q3b/OC7pxICdu2ntByMQm2IuIHkZoDNF4FwC88RML5GQnFbVtpyeeBR3x7lDW7Cra1z/vrU+
P+NREBwJegZpdtYkAP2LXFIeEaIgydi91vrDRX50q7/EOP4klyw+GjSw1AwMWtjlghmE6iv/Qq7s
i11J21MuXO8a2aXAsxj5DNneDWaJ3FxL1uGxMvkxQBQkqxDLYf2i+ftxRP//BuDrgVRvA+cDxSvS
aelUznJeZzvdZ/TWEh5QjSLCBnqjSenrfm4Omz3NGgbqb4LaAOVpDxf3rH1B3IBuTWvJbV9o9bts
K7PQmEXUlJ7fyeszHfdPljwlrklcZWAU/ujOPhX9wDLPGIoRY1gpV2GhSavA1vzJol68e0SBaqKP
lcfD7fQgJ8TvQW+g8c8ujPNu1wnXNsfbPbK0pCWi0BHyZ+rWWqMbxjq79yT8JqpUWGnqb1y9Uynx
lX4Ld6JdgkKjWPqShudpSfyOWJ5CjE+kQJwDWW3a/wHPvp2zBCpAiLaojnHQfwz+09Q11ZQ1V48a
6Cf8tZk2hzkNhQxJW09r7QjY803Zy8ixOuJmoc8NTUp2qwNEOhTMJiZ1VxmWfq9aGwdquVIIoB9N
L34X5NqkX5wR1toyMsliIzBPVtyq3F6Rbft7eNs7f+yDIn84OIrFU70lgvVZljq9zgbM0m1MdDrH
nfRr2wEvxzJL3TD2PYrccv7ezFJc+6KwJuRY7+h+QVyVqdrf8JiMnr9tNs3Ta598YA/sprjoJQOr
ZkEUoc3KItF82ZTF9vK/2faPukYocl6quXs8zuIXTDW6EriO3sJw+PaQ7jpoU28Iltc50Q9aRwtY
vAf4f5gEWx5HrSlQlyLHqU7p4iXB7/dDI8b0y7iu4Cdxt/x3X+huP2jLZtzjH1a5HmiWdtZSPVO4
8bUFaqKz3BUJwmu9N3BYYIUC9VYrcOgNlHZkxKayCCmjssBsJmlKwxjYiKQpkpC7fFWEcV8VxtkZ
VqgVsfxDsuGuRIe9nZ+mK+ne1X203GFWa493o6l6UTLJZzVMvGjQTi77014xiYvb9Qq0cd/6nDRf
4ZDleb3pyAQbXDlBGYZG9iAxyZKbler/ko+44GeqbZAyV5NFQP/wiAjVUgpPt0TrqVFO49RGQxMn
cjkl6JizFKxYMJDi4t7ADOqHku9SPXjYGT/CCVkQ2YC9Ix4r3xo2Nxgnfmfhh3WLAMXxTwhSdKnL
tNELbQmBFG4usMsUIsrWAWBchyUxHqgIBx7F4Hsxj7/OvSA2LyV9F5ljzJKYwNJxdyK5Pp1aWSef
8gIpB77VaIr30hs+A6dRZ0PP7uM9v1rYT4fIqYJ8wYYY7Jcy0A3tyWhyJIuERxoM5wDFJzThXk2C
q5pqeZMcahYX171peecMENXRhsAgne92agZk3BLRiiBA6dc5HCoLimQegj9n2aiotTHBnxeJ7dqQ
R4Lqrm12xPON1AaWU8vTcmKHQA/EB+Vd4aR8ajNWUMKZdOHoVc1aHckUNcuEsA91BqCKmTrj2UUA
etkqRnM/wlOrn96Ouh8f6XeRLPw7cfv3S2LjhIA4n5m5L+fnHdAHQyC0tV8I5c12Tm5+Usnkf/4l
R3qIMMu2mjBfOyww1WW4tNNiElp5DNz8VoiqKpuPUBOBVQGyKwn8ovhhgxej3S1GY65QQRqcfwAF
4t5YAZR2NCsBHaV4mU4/OvPgXi/kk9ABqm+T1NXdDcjTplefM66cqunpVDL3YSR0as7Mx7z8SES/
agz3PeTcDR4NEgSTDp5gsgxmI6dpRdeMRWRUfv/7xPKf76yd1oi0SPmwxI+H8tmZGp/6ngWbr36N
tgs2Z04Fk/wmymDy9sHbYTAz123bAEo8TYPOA2wxTs8BQI2XKEEJW94h4N8Wl1D4JxIfZ6A3unuu
dyvN120Q/LqNZfJ8fVhbmpov32RujYgKXoe6gVQ/IDhD0H9usGb+/piafxkAKDCyAzkCe9MFYOBW
J1p7Cu3DOrvYTmszFvJYnf/XRZ7a61JWI2PbdXhFAfI5NObfSNltzJNfioyIItFhlhn7JAxXtqyV
WmxECr63UJG0f9MOQFIWFTljw0Pty+PiNlYjcchZuYKWccwqihlV0C8n5MTOoyoxMCg+FSGsbj1J
KVj9/ujcjdglXbWkyFhNf/5C78J06KAZEAcqGWXUU4tQ58PzLsOlW1VN9dDgk3XwS/Z0VLBH8T+B
AASyWvTc9UFhAVeP0JSysHLjnUsYsAJVAyhin4WWe2zBhVWkOABVDx0AyAeTpxFt2zS52rGjyS2l
HTmn++WxKis1r259Gh2vxtykho81+zS85zwMLC+8ciBDYTJljNec5uJdSn3i+Rixao088Gy9X8iz
HvnJ9urYW4B+Nso5Da38/M1nHmmRup9PvSTezzSkFAuD2wnB6lqg7nTwaD112lEGomybWmngJVf+
8di4IX8SmsE+GsX7w8q0aAAETIUNd20E8RQ/T8EU6rRImF1QW4pf5iv+A8UJBHEMue4oOCF6XVm8
Ik5DQxQQfQHpLeRGrKStGQYc5ifMUnT0rSEu+MjHP3dEtbxXmeHmx7K+Hkteu1eW+ZrZzmiptCO0
vc6IuepK9oCkbP+SC4xGT9VOMLeAoKyng8h7BGCqD+S4jX2XxdZUXSA4Sao2xO2gZIBAl3gSnOWm
atnIWG8oEJyGeLtd3A053A2zzATAn2d0xv12/9lJxjAn3wGJTrLgigqqc+s2ng4gXHmCeFGdZ1e5
xEc9BDRhRsbZxnFHoSB+kJuwAUNdjO874RSVWC/8gIVqtxBuTPnhFu41pN/BK7nR7ePCArb2nDAl
E2KkAxibQ+3PnEVJzV7pxvnSLBNR3fuk6lcp7p4C+DIKublj1revpFShRVvsWMZttIXj8+yALtO6
sepvM9STl2s5YVUwEUKo4iCXREEsP0CHbEMO+UlWBCiEoT+x1APDM63MRC18EPXHj30SfL1WgMo3
KTjJhG9uh052KCCt3uYD+joja2lXTGc5GtGN0jsComH8eWd3wlFIqAIEwvUBbbx2VwfjcTXRiRa1
QNGf/AQR19Ow+eR29BgRPoGVS9w+Jj4m+ZdhFh/5fLSBRLje4JIW2nACU2bMgZ92dWA1WLbg/8T7
xXzrlEtIhrWaknuMwxE5jd7IPIii6ey7Alp30Wc1NAEZVb5nWeg/QHopKxjqwziCcD9e0k0beuXw
I/+h9ttOsX0LVmxXRAqR2VFPtP6+R4yzqO94bm5Nvd9LI2ugsa+kWH12952blV0GOQoDSF/pWsXz
WwdzoXNw9BJ4xrs6Ih8LU8CWKZH16A6gNdPA7SMUP1mTHOQgfA0f88hFGjSy8qT9d7RcHwDFns/P
buCyTOFlWuQQRNZOfwTotdy57gUzA5Xq7Vq4vB3PC+HTmCRDmH/Nt7VgA7qkDIH+plndOp2UBB0m
c2RWzvjPZ/mm5okRJkONMYBOyULMv9twiPY4hz6hUkFFqDoAxRbF3M4104N7mzTHA6T0kUMRjVZN
PLYOB9xqxwSQ5FyiH3t9NNY7gQ5FTQryHpUUL6HLB5aU7t9wTSCX26NtNJ4kcEL/3xv2Lvrz1Vm3
UCcDhiGcS9EKBJtdiziMx4fcKk8ObDIxmyP/sIK7NpsjcpusqhGPwOTWv7TZwFlQIQ0AzLmljVdC
oVh5xJb1ikDNxaEW6JBEazcgFN8YHA1CzpA9ietOI3I7zXOgoihGc0tgFAIoKscmNY7SwnmCwxLp
Ghok0w97I1/s2wLdnyViT19blMglLJvB5NBFL4Z4PABgNxeXjICRz3GwBX/fPF9GVkHBuI+GZYlt
HxxyyKPJTAIBn+XcO1b6gwYFeeHnAJawomuDQHwW7VcqD+NNSLHh52PahJjwzfKNZFXg1mt0SmHo
a1lws64X0mH4R6IwpD4MtfwS84QIYRhmSvn4cjDWPrYrjQi96lElwQNJE4+SRmU1lJysp8hrpjU0
zg8/UvN5rQArDJ/t0NG5VfBltHS4s/l81XJj9XlphAP/rW0RgaNCxd+nK71TG1hgOWDbUaLRBEA0
DcQOZW1E74QCLPjDRkF051O74CZjTKusdPcCWZDHfIcnUIGW5UF0/I7OIZh4CX8UyAuxo0T4r8Lc
ztKuLzEuHhw798f8nhUNmgye/fNTHATI1LSuW2/InahK33dTfOg+r/1hbTyMpcsyaTgPOhqwpMPQ
5XSdEFlPt1BQUYy85GijDomvjonTBkKc68OC9q2D5JhVStF2fknX2yhOQ5rGPxN681MA657D2weH
V8vKIEqchZwsmKnPED/41a+p5vqmfHSiDjcc8qIcKTpRWrlGFzS38J2/fo0DTaMDOUpBfPuz8ieE
7LLUhknayWl5/z6CeewOSznBfsSb1prmaohhIKQYlKmH9N/AlospEzyYOyWIcPiZg5WuH1aeVlOL
Nsl99M7kVzM5UuHp2vAjZDbQrRgOdCH/lRVME682Ang3v5oAGrvKKwEzUsaN1UbSJqDv5EXUtjtS
391jJHymrWA0xunf9A8Y7GUcwt4f62/wiTIPPmKEX+EQ2UrQHzPLeAInu6raFRzpmgARCfkAjp0t
oPOnsEil+SwKhqSQvG/J6LIoR9wu/OAXgDvZxwrBalGxdMngSHdz9wtDRBGGhQhwoVGFSYrMuxlH
7k0oynrCEN33T7EBoUkNOIvvc6cPRf+5261ySucex7aELX3vQMKqgtV8j7yQn7rZQR5tyfA4wbKg
UugIRmsm+VnTwR55V2n33iT7BVzgNWAxmtRMCfrk4csqm+I4qEh4aZTZ+cdhzUXgEI/G6nVPgGR9
y95pxsUByR+WeO7xymp7fbYsu/YX4qwGEinU8FW7l2bYZvjj/R+De8sFXPdK4is6b4oPFeoancnC
7LgjIN8XuFkmU5BZAnKi23vIp6lC/SiWmIF4eQm+Th/KzJFBAaaGGZmjRDgJnnu7xwlSO0v6Acy8
XjETeziZjxzs8yntBTLN8ugATqfVWg4fiah+uR7Wv76wq2qCuBEtkBQr/fBln4uff6FFICsDIahm
kXa+UYnrTPyxcC+rIPhWWtf4emssgZkQ6o2K3hpzLhQH42hfXuM+VKrlOrsAVPw9q/m93UxW88KV
S+4vVJVH5npbDhd0Uyy1S5uTINmh1GMgsxjnsSWYHJjNMqUbfnSGQutwJVmjYKEoV9ZEL5dXgG12
t4Ri9ta1UwUomeJhmTm3Sw+X08yHW05zZaFj+hgGNHnKcKt38TfepWyAwwgGwZbi4trV3jsGBP4W
ELTbd6xg/NrRoz7M4z6eHD4mpDdk7tsq4GoJoihWCFlOiFwQodO9CO1gP3o8C/rMJvrmR5Cpxicw
HgNJF0G0J9Izf7PmGemrLX8RoOk1HQLLHENAXFkZOUNkHnytN0oWMKCjWiKiJ08/Pk+WJe1VVLr+
5KdkuKCeB2n0J0nU9loaRedV9nVwSJiQ/8fN9dLdRUOOrgo5DaqAghZYigCshgmOzDkqT1Jw3bWK
iAC52uXKd6nZAzNbYnpdp4GwkQzwtux+0MtcMGPNMk1D8xpM49iPItQA4ycG3HUSxyPqpLgJ8w5E
+Kf0JVYRYzozAfHYj0u9v3KSmw2rQ7l81tj0ZhW5Wg/O7jQ9Xvr/wFSWE/ZxKoX2xLQRVmOsZ7Ap
yqao9ZWpFRucOIjVaRP/FPok1X5qfD97wkN4CwKqj74CQF8MX4U61CLbfISWKFOHABmm40WZh/xm
2LzaO57BQ5+QFhcR1ntq3XCMROsGZxZBWNHnE7Lq7C+/I3+s3gyKbrDg1vjHb3VWs2XsI4oVzbvy
W36jBKu5Bza7Uft1ZiWF3y4VIqXUux2RbBoyx0ovt1T8dsTu8iWOkDVG1O8ZmUf7NQZJL3M17+e+
Di5jAZIdSZswAIxIuVHtxMWuuWFdfyeIKsg9VcZ25n4ovuk2m0Pk3mWhRKpTisT7NFvZMDsT/und
+BhYeajPXa6MWc1AEODVE/Vsyn0CQoTQkg+gaZbXBAHAKDFJeYGCmgj+4JX3D7NlRZLnyI0gRxND
Xa9Z6VTsli94xfgVorr/woeFemALhRnNbPpY4T9pI9fW4dvHd7wz09AUfrAIbEGpFdhS/GVXRa+N
TZV+B7ez8M3Pg4UaC4mRk0kuTWJ04qNBTZcRbVLEb68QS45ThDJLI/hbk9hgmqjZeK7Vzkt5IaQ3
pZjcz7o8imwLqlbBGVI22lck5AZTWmp5qXANPwltob5q74MBnYOn5MlF8eai7odVOvy0SdAQJscX
HRsDDX/lKz6InhSJzcjuypz+IMLHcSGUlCkcuuTRn1LD4Pd7a48GsG0zA6zr1kgVap2nyhOPP+uQ
xfy/3Dn/p3miuHgbmfBW8/EubOgL6q3va0ythhcNuF0Uw1vs3QdymSPbvQK5fU2f1JY9ARq6vsf+
qMDnZExGE8xIVTQssFn3TSsm+u872qGPOFqZae8ZQNz0gLGnpAVugGoUowh/kVY+ja8pbeiUeyZa
/kKVke4oti0Rj6BJyTbrMSAhf/RrwsUo/qMhTwLGzFwXuD56a3HvU4oACp0BmzPJtJbWONMXFcps
1pwOiB1yh4zljlgz3BedDyyYjZnHc8W2nCZqwK3Hxrrxs0XtxIpFMUxsfGiJl2BDVFfRo87QCl+n
ZIcRnqPx+d3i4wM9uXALY7Jp8SbhCna2iAUgsZp07AgIZ9Zz++pt1CW9AZkdihQ7o3/wHr2eHwaz
ndgROrVt1bLMLfGOiGjWUb7dM+mTc9gEGtiyHEoo9Chh/TxEwSkG70YJ5EJwh64rBFZqR2is81pA
5mFFBlVRHySYekWwjby0VPlP2M79pF18RAmfpx2BgQdTi6qW4CGP4kLOnvritmLD0o/GUUgm+/hP
NdewCgL/fIJdjyxIQb91Z6gJ6BSvOoO7tLviS4PkS+MBlwChXaJGECKNCiD1V/0P4MWHZI4p18IT
3CFe0g3fH1RI2eySyH+Ah19nI0oad3YDYoBx+cQ4Fz1aS0a4aEMjmBR7rgvPJLNaBsNTyLKJ7/Yj
PqYig1Q1TRCm87AfpZSbyjfE01wT2Lu/h6qlC0oxDPKN33wSy0atgszvc4CiHq+gY9eiBKDUpv9c
/vB2roxOCxyZgYnmvVP0oPWlyhKswUBTZdLvoqZEx1/GpiHHdzrdG+UN3nSIbeYknNxhDuMyUU0Y
7cfjT1h82QZo/lq7canwaqMV+aGnDmRfa0XLuECw5yRPzOtc6g5VkVlFGI+w5E5zuCpRnXDKLKcH
4w0BjKgi0lXPjLruzBG72ZlR8Ki3sxJO5NIlUn0GMct9qgA8kxbB0WjBE/KJS//bNHlPJvOOLL/b
9fSSYBW7TgkOT897iUtOPETg3U+1+pBJu1HWYQh+IJidHSw76teUAdNtpI8xYKdr4kC1J3MPhZqt
GIE7NV0bEWyg0UfxgAlO9RfNFKcCgeM+kqvOivKqxKhNt/rs2I5lODKVQ8xV/C0H9VnxW3tL2EmA
eMp8t6r80KWZ1snRH8vs/bFWRu+Ld6wFk6d37b1cfK2OXLt7mRHZJ2SZQik7Q7/Zs7JtEA96Q1e1
QYYHj465QPep1HQDQE47kyd7SsRHm6vHVnOB6TTfLFPWirXAFeDPuttRlTMsUbT280YR8jan/QFx
dK3gxCJmSL5EbNVzkm20Sj949lKAC8bVMAvgOH8ktqrBbsQXkINg6MuDOcAyU+0s4GfURw1jWXgr
FYY/BH+1OhRDskcLlgS9gtVKoPWf3D7ReDOBCI+jKv1/v2pGa/7WVN9f4gBHs5QfaoGtRLBaMxRI
jf/MINifJtFG7EmNfcsUZuAW/PJsQVyRtB0fQk3+OHG6fO4lryj/lTsT/GL6FAE+v6Bh0yqzV5nC
e8d63lkD/6QB2vrwiiXr/CP3PxrzTngBj5SrBSIy3i3xO/DbNTceaLtCGdG0Vco+FvUg248jUxtp
WB7OTnW9SKGfytOS2qV9N3bgDa+LoiYHXEgh7OKjhKg3+t0mzIGKoy28PvJy+IkAEYpwJaaMZ+ff
mYce2G++oqgM5gI2aLjOOy8l2JVc0gFTTzO2Gof2sbYqmN2YFgDxf8T0mQKWEP8KSy2B2faVC5sc
0/O3Kx9R+BOBnC41sPuKgV58qFAT5SfR7hlIBbBTCPJ2A1VurN4J0gDXeXA9WhjGh3xLmayKEldU
uN5bSdpKpswHHwVEVcbpbAveA3U01ShQzOypWGEUo/L3o5Iav7Layb9tWy78N2d7y7FSCbz1kDKF
Jz3E5dZVhesJRUQtGhTzXMuXMTx+xTszoOgB4jTnV3xfJbRI3VXwu3x37ff5SMHgNPUVgpg6XbPv
H515hPrfUAoyYxC2yaE/Nly3HJDjbQf/Ixna8YX+iGwYlDBOMhxg8Ovf1DxtWMRt9HLaALq6DBv0
azvwdTX5zu5iYjXY/j2L31YZYrKbbsRv4Z5zXW7dtTzGe5cYwUw4ckKSwxX8+ZoeEOg9j3un6pH2
WdgVAaDDw6e/fB/WnOzSglhrTu54mHNz57mLzcqL39jJLAKOiLAusqsxcZwYnhnJ5134hBsG6WKT
enQU+LW+WX6IRsG/9BS1ZSiae7cD9v3KnGpFYtNbVmBx26YDWxK2P3DjC5Jw5GeV2hPKEPQpdHOF
kDQh47trHxUFpshX4PLK7gTHspLwChLfEpTrky9vz9yK/8WT9CpeYABv8Taw+6jm3Exk2GZpX3xI
jcTpzIQ/8nyGFzhZXNeReUr7XJwjiVJK+MPde3FcughBQNO4k4TlRNjeKXUbQBXWm3bIBejoFxzu
4odDaX3iAqnrWkDBIYDlHYZYesZwgBL+HYJ5uR5kpr+DU87PTtANPc4mh88ALBdGsII3kYXtbIyq
Hr2NMVjCixUQtLG99yxDh5GWtSQkQZspjBQguYRAQ4nRRNYRB3okOuEg2CNpOxDL0louHtYShDKk
+Hd99ahMwNMP1yKrL21pGQY5Fdyk4jHnllfng/YZYp9G7VvzvgGbrdzjk3l8+PlL/1QwWCY4c/jB
qvq8/MI70fUGU/GPkI2DM8VdaMJHwKzmEGJ6gMRtLFZxC6vAkqq9dJFXfe/Cpt0pBnTzSbbDiCZE
/UWg/uREXsuZ6EsP3KCUk6GxznyIfDG/4td36qMABxlZAKRtk5SUAxMfDkuG1sBqqbrDABs5XZVD
VZE/Jk7OoWeCgdZwaYBpVdCE2jxP0JqMfryLCigH/ZeKJUW2VFW8OlozsYQ5oIt5m/9QdVzLZZXM
EUZBdzOzKT/Je/Zd+kp/1WZaC/oA1cGjQQ/kaQQriXS6xcPJf6bsnmtwJibEoj6xmw6OAIeoNF+w
eL7jR969tURry4O5iCoS2uEwGsTixpGWc/q17nElvCB3n6CunA8+kLhKhXkky/95z1XT8FaPcc7Q
jm2a/jJ9qDuNFErzGdlkFugk/iCfmtNxesWhe5XiV7qSRX9stapCkPqbehdVgsY2p86EiV794rc2
N6IKaY0fEA05Be2Va1ISDKcU0B86+IYBsFzZ10ZBz0tEXX5PUXrVw2o6wqYzVAEMckMWfgrgzgk3
D+S3Ly1eJ3U3M4FNZN6lPmTEE3Y0sr4YyH8QMVslc07nD7VQSwVFbUpvx2UbbS1tNc7wkOnQ6KYA
u71iMiFPy2uv0MwwPWzhbKx3McPen0S0dc5715f5GUgbbKfFdB+aWXjOwsvkiCONTAbjq8E6EywM
3ZV6ycK5YvCRIMxlb6rtx2DmxEYnFY41A5EraYxYbpXqDQ9C5i62YvXJ2aeKDGgpqwZc1+JJJV9Z
2DZXUBg35Udo4gJ7DUPRxKJ08E3yTt9f2NlDhNi2G+u83HXXuc5mOU+9+Hd4PtScBgPeJAl0ckQq
VbC0/emlrdVBRbBFM5SmLyvzN7uLQS5ltAorU6EiwnJkKN64qQMcXuziJAh7imhIb3/8Y4NLRwhG
Kncfp3Ee05JOZTpg3abt+LjLpE3zAaA8ThdR1xaziNMJe0EmbqaTnsNaE/WBtyX5+7A2sdlX7x00
sfx1Tz7XAh3My3x0bhWJ+0IvdV5U2n2G7n5OiDwi5CvZ3WW5kyuxJ5wDK+Mz75RUaWYKRi8KL8RD
haQaJ0YdSHM552NShAXuQoVUiDOiYzo42Uz68Y3N0+wkiqa7xjSHfjzMN9XTSaodemQ6/DvKI39s
At8mKhn8Nlp2NJv4zikmkG6AHMDUBnqsNhfrstEEC/cB0PbswfEANkgRogVrBnJXxiDOYpGlwuz0
op5sT6Tc0StiTPFt/VUEoLH8+pU4X6MBtAKcFvcIQvjnoOGL034FjJ/X27KT9Zw6iYjpxwAxeold
3SCowfKiTmleFde12k5iRpOdBABzzDGN7CaH5CD4kH87AhFnUg0MHlPBmNOsgLMSrNEdrsPX/1Eh
zMoZgQx0Bsfnubc3Rx1R1m8c2Z14F/Ll0TN0Fy0aeeSHyVCZfVCp9MR3ueADwvezejtbErDCeaEM
Pw1WbRBFdNKwylaIUCWbYTYHEQBTdvOF5fxZ4e5WdR7TdQ9SFwJOpXhnebvHG6RaoXasUBQqDmUy
MZiYRUSMrJrYBKXzwYVe6iAF1IAiT2oGkj3ot2LL9LLqvNVAZtp/sXCV5Arj327jdTe+JqS2ytG2
6qLVdeXD8kgU03K5yAgke0AlbDrDkKbONFJyhnbfehvPQSTze4KMPXRTgRtQqYPpFl17UmdKlbZV
+VexdynBja4Q2o90+393pl8B2d3AwK0jptkJ2lO1tvda6/AclDwiaikN3k0Cm3LwbaP9kwsIEZG7
vbEvZ+vVp+1C3xR96ZF9twDMS2YUUQhE39f0CmEbua2CpeXBnX3G9Sg1aaSAEky65ovKFJjMSUmX
ySfoCRGhj67UG5rPqMVwl/dmsaH1pCzgLrhpxvUwp8nb/MhOS2rBc1hwKmlZDJcJpx8uxOs2Nf0u
7FBZpyTMGLjCVcEPU2YUB77GiNLzib5ngFZ1jJrZ3bvKQSIzs3JmWF6+T9yIx4M3nae8C9UZjnyI
Kea+UARnSRrIAO0F0Oy3TsQB1pe33sGzbXupOgYr3byvWIk6ZqcWoh0CDrSIJdkgViLydjyHhWCQ
c4aJLPldGfDlYuWX4pCUsk+82PKvvkJCe2feXC3cUNgiEJr4DnRjIjD+RGAIJ0d5TMTfS5vkV4RQ
xC0noPUPR9A1oh9Csl3zxJHpt3GzyT95HczTxIumfGAH5EhmsB3ox1NrUmsHBDqGUq9efBhmOA08
Cx4OpsIe8iLEKcw1gG86GbRZEGVDSTnoSsjfTaNvY4RioGKzZqHJGlUKvD/awltB4+nwHfQDmATJ
8F5ybRuBEeD3ku9HJg79f3S1pbDrkGfcbwnm8vkDReKLTljj7pc1a+iV57vkgxkEzO6Nts+AQcBZ
sibZMn0anAgNZVqB+dTIX18Ce4+oEQdFklLrsnq0CVZszhlsStdfuRm9nGoninfx7mSVj0F5xsDj
n7t2WFIO9zyBVLdIpe9ZdtwDvwv/LiqnVensOs8V+mXEsf5jBjY5vYdi88peIKuLRLRaefisRivE
PeZokLXVSFYCHQGLHeyoPfX9Dieyq7dk+wczvYGTVeqzT5x6NqMAY8B6oPNSugQdieg1qk6H8ww5
qZs5GmOx3wRcSZya9E4Iu22kWd9IL3k304I6DQ/rYme5clmSnYrhtcPyDpF9IQp5HyCxMvpn7KtE
kdjXBzX5qFZvaMeKBSq5qraOHyCv8pjyrl8BljTBaRFZ+4cZvLB9FV5WyHRmA45XY+7ccnhmM6cp
fnsOvcEkhWzMazc+6ZBa9CTFhHpxvkRO9tXwbOJd9cvmu0uC/H7oY0OOEvhIcKqFwXHcar0kggfr
vxUDqpozMFlgzhKbb9kwAl3sbS/32kdYH/vh5yRKL45aePFKTGlHpCuMlMjilc3Ntyc9yKOASU+o
Xw8ImEhwNutggCmYaw3lscFSpK+Yx/wXMKSDlhSLqQ41w3Y2m9IFU/MVLq/DMyAicB/Z9pU1eZh3
93bY9P+Odx2+lwQCCaV914ljBcSE8HmSyV9sBZqbeUtfFCP+NPDYK7M54XnOs8WoUieh12ZiqNNw
sFbXa65BBEaynpaNCXxN2wuLM0xQynjpz9I0D8Ds5CPwgf+KCTX1A2nQCdLx2nmeAd8fhJFb6eZQ
L11+TenkO2sViU/LU36UU/NAf65NTXFzeaTY6p7mU7FAb2Yh89ItOsShHIRQzWh3AGwDxFbwrn2u
C9uVLd7KxBmctmFi8GjFC2sUMoiFzGDZah25zjBlxZmMI1bCTE/i0iExuMjWHwOH0RfHH3uM2L2L
yBQ30asm/nu/GsJScLvA0TjqWPfXAi+wv4hIz+F4eu7hIy1qa4YKUNyIC6Bo9Uaxv0TxCkkp8jtA
Q+m6lXgyNm2JGfBYTTiWVCcZejS0nlA+fT9zj/quGbpuaEjY1Ac0I+hzi/hK1x7ZP1mizs9WGbGs
prr417t+7VHquOWIW0Czqp6mjGxZrGOgf9gdQ3DaeJMzKESEzVQtdId5l94hX6k3JN4yI0z2DYP2
pYDIxTrFHc044YvSCvSI/Xz6tNrNaFb3KgdICUcFR++KlsglrWAzotMiODcH0ikb0tGoZP0vUrjh
PFCQhzabiE6glBz3eSVG82srSiJGXDq92jRhskDCm6S7o5PSSTZZEfm2N9Ew5u6F1QZN8XANreA3
G8z/fxrY3YLk1Ahq3AaSyWX+wxyiEXrEHHUHNWI1pEH/Nv3NtajTUlaDqEox5LVOca/R3INQJHfP
gdf9Uik8X66EXTnmXzXdjq8xkc8eBaBznG2WuQIIkDNbI5EMMcKO4Q1nH7vdhJSkzKuL9BSqQTlO
X+X/B934ng1JmQKNXPulnB+QDoyywzZthfixZRGk3TARlZWB+fxbY5scZdGkAm2cH1pL4yabddDf
HoL0N66NG/qEAUVNxMpFSDob4DpLPywPVHFBW+jylRKoRpAYqRZqoRmDQXgx7Ls6yiCoiUnNKHLQ
r17DFc8Nh7lgv0RuvFwy1iTZk8q8zAdvTPpfD5VJZD6cN0EccTR3YKLOAF7lDZi+2BX07LHTNhSz
grFRLGWtwdq62dRNxPcbjQINZil9YfuJv21JRJDj6yPM5UmSQPIx2EpCYAwB8eF2hNyXpsu51Goc
ul/jmV7uoTAY5PPBs9AWirXF/QIKZRSSHMseZhwnaUEVrVBk14iUgr47YCyF07+hft/bDZCA/xdt
KW+MlQAJKdcxAy7SPu/hzU1ZVset5UIIj/ggXw7EUDH1AlZl2MAfB2nFSgSeG5SQDMohPtPqMevT
UuTFmWiVumgF6gmLqtiw6cdnEfTxwe1OqylyANB7n49EmYIth+LD4nua83amv1f/1FKNtpbmZ4Ei
Sd2ZZr3v+n+uJqogyfJ782JBGTcQxM/TUYtyXNz98DND1JqiBqLxoqzuy4PAhE3O+v1EpwdpqJAa
XG0+eFsrHwHfoeAStE9CFDQYYzQkmSN+mACJ/KFy3w8EyfQlm06Tl+MlvW+Oi7nWp1pGY3bWvkuP
OKV6N+hUk+6c3milgRzBVTSvutVcKkvjnDWNVm7bdioh1IsyvEasUkf9MaDC1Ct9FjAP6hai8MLd
fwggFTezXapWVcRUQBvunzopkRogl47e/Gu+4DoObO9kU3Zm8ZM+8xiol6DY6O7g85Uye2OxkiAG
J6MxUX064XxjjPJaZErvZmd5dqT4FIzvtIHsXivh5QnD2KrdiUIomLvFH8ch9kfzWKbpvyK/WLrd
Fk7AfaeZa5TU9bXJ+NzHKUNm//YP5Qqb23jMEvm6LoHAhL7O2ic/FLk8h+/fvIDOljOpi/BwdA4Z
UP9wwSSSmp3QDmeaFJZBY2Lr4ezxeg8/1PekWAPNgzq4P/pLUjjbEW13HG6Yvtl61yg4N1SlqVu0
8vQUj1fZYgfaDhbB8xzee/nwR5Rz4pD1ul3TLvXQSN+5MzajPM+Am5SgOUHVcTaoLGYGco47pp7E
zKtMlfxTwsrUDP+rfWw+gieUdSIkhPuR69oWXdvCZNkuwxFZw4tywpZgv6sESKFi0qiyGqPc59+E
1OAkarezHx7NVkqs0VU71CpXYjctfWn23QNly/EjacfsIUfGFktOT9dM1eAcqNh0ipyXPBU7zsKR
srhW+pgM9E8gxtA39KRhxs3ugCKSeLScDa45tOsKfEdX8nPTMBsELlUQuCGj17sBRPHx4524SzOx
Til+m9dxZuCAXBhLtLrHbsVdQdtvXfRsF6UNzxE4nUW8mE2PsBk9eRXHDGjfd1cDH24wTOz8PMOM
v5zlvFL2lOnAu1alKy+5Jx8fRDiQD7L2xxFfV5xvFzcxuZTnUezGbiBTJTH/iQjkfBtAEJypLCZA
D5AEZll+Qw5FTzL1rxZG6HxYe9k2SImt8ejaeAqVtIm2HwyTjOhAbHEW93AzJwkzBM7WVq4OqSgb
vmAKXGc6MAEmzDAQjRN87iW9RJREv9jLAeZnw3bo9Ohh74FTSkX8mcz8FzBlL/x/31waNkpJOKpe
XXKPz/qbYq5cYMGFas4YkrOWUdYuKh+wRlJ9XV7Rxrn6HBQNTwGL6OrgqzuLAbImEArRJzALiSo4
eZZZQ3ECagzSu9bUwSwiyGHCVQcJqEiZaNd4tgPMli97DFcCCAYFJtIlzVS6o8EA/fLUk4ubZKA7
MycmGez7ZwE0PGuWthBkAlfMhL4WZ2W03h8/qtjXyKC4Ao3L5N7flp1qgYs3Cl04a6Ug0Nd+OoHp
O9P9U214yyPd+i0L9qs3g9Z0APDrXhhnnUAe4+VZKqctnuH5uiSQg1XgsiDtV8oTpWK9IcYULE4j
SBbKFqZqlVvbpCBO76inbgAZLyzllMokuR1L3WwvY5J8IvFsNNk2XsmgcC+Sb0MDa62iTDI27iaL
P4mlf8TgmXytjPxRKKEjaxOkWUa+amShSHHJ4Yhwg83D+119FVrm6U4oJ7VhUALoprTmiPF5nMLJ
MhqzJClsm4FEzB0/9UlhnaQIycBEMtB4k6fkkgeQp6QONfz5b+CN34FKY73YpBfeV6dZ6p5H6fed
fJIq0t4E7L1A90gD/iv2BzoJAsSmPXYrMInaT3b8A1GkfAh1mQhLrnOYoZ+67j+eQY8a4J5ILQPP
m0pib6sn5B3IpyzCEekux/tYEjRh+oHqOQ355amNaNFqL4WG2EOXFVHa4ozB4iOphK7md5BZ+hvg
3jZCRRLBR+koTkL17tGpSPMiIKh8RR+KDWQmh74OGWXUfjATc/r3dqTqJ6JkdbkFsfGrOfs5XaLQ
7VYpNkwdU1utfvmKnJJ8v9wjqoJjRl4yo1WS3Bi85OOK8AsIsokfNwBVzAUt7YLXsS4S/w5AQlBd
fhiZZg7/XVk/jHEQrMCBa+U51lH96S/brjN9+4I7zcSowlmP10WnogADSzeJ7gma5MUwuW3ac41i
SNxanmCIzzXD0VCkgCV8buowXIrpjluaIp43LkN0cw/OQzFu1ZoVD25cJEaf/zJnFzvyIvj8kM0r
xtsxQFTDfIfSDeZG7dPf+8a5QupMNxvSq6RMM9KwTQPp8fTWQXYUJx/9mcUatUl06GIAzEllnkdX
jf5dYduofvvzhlxZPEOCDx12mJwkn5PtJQalXcEPegExJOhwOEL0F+AN+maLkb8Rk09oA0rdxqB7
/24dVzmYxL9BnPy87xlmhqvGCygaUBQPNtZH2SXlhGwbApVVPoxHYSA/eKYYLN5dKUekikzGzY91
sF0Daxp+y4ThTFR9c4pWXCXsP0EjALn3kYr9fiO5RotwrqSeAUa64DK9D7Umi6Gp5rODN1m7dT//
Xvm5ib353rmIA4mbNbKrvy5yVDmZSOlGzZ6sh3WTGdeFNwgGadcikpT2gjOxSl/M5DP6+wC5l4ic
kylewWD4I0jDwxP5NJCIkPJGsVmsoA6T7eJKUPM0gIl8kh9zMGqqE0HGUBp2IYy+rXplL3I6szYH
b1rwUo9DbZieawAtaVKyALPg4/M6FqXd/ilVaVqBrmNs42T2HNkOweD8Gi1p0xKKdtC3Llzrvte1
7hw+Kwi1epOTZtOrGTqA9QftATi3ZSoAHlIz/WT30kTL1FLOwV7CY3geWryYoA1aUK1EQdg37sJm
tf9NxGrT2W2yJUWVDnICZu8DLds462uS3RdUuVocklURekCifyqedDjYBQlq2fDBgLgnn4R736Ez
SHmWNXVX+BteCuaEb0H6nD7op1bnRSKzHvsHwAeQfLOhGkGCLauNk9y50UzSmSGUS3S7oSmaQwLa
Rrm7ieb4uYbiQsz+K56Rq2lJjTdovXprESgmBerCL3gItSLw+0xIfL5LFnB4DVUdgMKSTfYuCPQH
wjoovvzcKucWZtLnGOmR9Anr5f3om5yy6lRGAf4HlPnC7Xxu6bDWotRxIJPXnw3WrvD01PftqNjW
JTI5yZov2LM4WubHDnQ9830e8O8x+orUzWSU1K2y7YXAnFb3AC2d1Ln/14DrFeRdAH7gxAY5nnWw
dFTSKbgboSWrKor6j8bliTza+tLQt+3zAyMZeSlA7uszymSoQQbLPtikoJ+bUqyOGh4pSQ+/ERT6
8Dx2aTmVYOMyC7GKLPTXm7B/jxSMAfc0KZX035ZvM4ULqryd6DHJcykTEtxBTv8WsP/F6UWkkIa8
P+41fmb1/CGhR0KjhUmVVydRuoGfIJ03kA4DEdLtNMMR2sd93JY3Ff5D2JYaB2hZjx8wYQSQre82
xoAcWqGLlZ8u0M+kvtBR3HAHQnKPO9tL1gjQzrZfdoui1BeRnVhc9oooFKAPxfFQSpEC8diU/9sU
seTiHEEnY4QORSRfDdKPDEC1fxQxn8h6gw1ciUWtQBKDsaqceyQr+AqLh79+kHaf7MORXr1Vvuw3
bGF51uHNOVL8biqgCNdryjonM0YD7I65cyFrMq4j4Z4lyjMTtTG/uQEjb8J9Rmb7TgbTo/w1TswI
VDf1ipY1QKFwsPeDuVji5fDdZjyf0MTErk1HTcaMU2MT+C6C7WDkymMzK9TSOBAxAIgf2dRUrkdi
i7XMi5BGeFlGoAIZ7VI4bnMY5pfqR0AIZCu+u606kUBgUNO0I0kAocY/O6TIw3DU67KSUlXOqKDu
kfO2Gbhj0YSTKb6HD9RhrQoqmtx+SXD+VVfx0ALe9psbaImilfnZsof3n/fwsTlpXIY44UKFmshp
CSnz2/MsVfr4x0PzDhGwWhRWNF6Auo0QNTSzRIuHxPe5XQQEJA6b+G/05hGhJ3EW7wV+BoaQjFM9
9pXq/oZQchxM9bF8068M3YVpATYQMUxq73dfHGy2PURRzcoEVJAgI9s8OvpLfa6Rt0bWA/D1m8Ja
cHOY7PnOO4+4hEttEXPkix2Jz+QvkDi/I2Z6pwMKxfz3jDBrIVv7hyC3sAywQ2qffVIubWUQabmV
/F0JFSvmLCoGaPAOQSh6ensRYk2ZZlr3FsaHCYq/IyfvQkAFtV64Ur+Geh/70hwlpFpmqNiHul4/
SAzvUTntAQdqWtzie2fiua0xavkhZ0JRnANBSumQzmqiUuBOJ3hB/O/RMp3hqu+tamKQ605HPtdK
E5dxtIArF5Aa6uJwBR5V6CojYSbpsIT7Z1ILam7Fr9sp0z/+hv5xrHClWQ36P1JrMSOUn3pOiNh3
KckS1CZ0u3Ba9sR1EdDNC2h9zCPzzDrOKzdE0qbQGHgqmSJ1g4XXMobiX1VS0hBmXpeX+VXj1RAG
7/2G0mNIlWI/yGEiFp3tmxE3UgSp6aWpXU5wH3jnDoP8sitVJnFLb8kL9hrqJ6HI1vM8qaS3K2al
oCro/I1KQ5AYDssWrooYOlgrYLR89RW8AM1v2B7D76JDvcW0P1KgeJKBTxhx6vz0gFF6vsBiJX/n
K1IoonBPdGlu4zv7MFqBtMTGNTlMzYdX5K4QUkOUX8VXQYYr9V9SmYJsiVVhJlrDQ5pgyDwb3Ris
0POL2pUUmBmQ0kW5ZH6lvcqhM+TK/gqN2HfbP06xw7vckot9g9SAqYSFgsVsL5TgsTqAR/2akxMc
b/CnOwJQPqgwHye+/ii26n4B0bt1IxZT/ORo9YfdhMqaJFW3C7aUnIDl9gpVRacA+4kX/v9Wg5Qa
nUmZCAARunuN0PYgDXqmz76kIOFi16TGkCTWKRmOKPxDSLdPIujkBAutx8B4CkEmKTG/MsYiSWxP
UwBBwEpD/SbUw0WJzY6dEonjZ3m7Ey5wyz/n0QYLlSbBrTvdbc8v8CSGy772HB8Uoy3DOtv7GVAq
pI5owdxeFEDxAtR00DG4sgke6zvpB0RBLNQIQU/aaI91uSWTXErKsN/TgnskRxqrfQN1o8VMgxkU
KiGzyYUxxDuKY9xcDJ7hYKVQaJTa1p/8+qPYVEzyuYvFwSoJOjZ1qO8vKz3qeq/xnVzDp6oLpPtc
+RrALlHefLSdNcDeslHuLnO1wUng5w3sfmC5VhGMpDL7DyJ+zhgWCJbw7pAdrLRx88si2NWlvxeS
mBLbXd/HlZpoNrBsoY+nW9SeJ8usf+f/53M7G3DYr2eHfgti/QJHa35BwAogfOrzRYMbMgENb1PT
QyBeBrro3yeJNUN5OGzo/ax6U7MmzmFpWzTZgy3/BoUDJskMamQS01Uj+jRRMn5HfWbxWcgF7z6H
28YlErAxQ6mAaa3pCZ0c+BalREKnjdgsDZceKkEBg1UZB/9hTHpE9kysm/esSSZplNeEl/gK28HV
WatfRSzpFKlICfntBPBmzSHg0cgbmk1zxxeyjP4FJ2ATbwuaTDopzg/kUOyOk9GYJJYEs4KvL2GQ
AJTKLeMD5VtwLi93+xzUEwH8WUwsvxMpN/s0wfG/IzUjXOHEnvZvz5/MBnUpTypivwSuLmBEwpv4
GICAmdP8tRiu2jNbxYUvQtusXCOSaOCHg9RakAFbJXqP2pUvNooShPbkX7dgPabFTvf/ZHLBRkFl
9Hah1hlfcB7oxVBKJrH/OlIjPVVLmj7AbqIG2hz+tD9vbtk2N2FtNIgPwP33h1B6BkKT0cdHnJ7F
rkalxGMTrWvEnjHn6e4ot87vaOYWGuEnrxms/1211ASTMf4/zB8Alrt7g/Jq3mXVadxT57dkvLh1
fj5F4IpCiewg5jOL3GSpr5fFQLyj9IjF4Idd5a2gmoPr8OodH5ksF4NA0e4SDoxjgwMnDkxr8Pxo
Tiv7RJbzI8y8rvAE2k03xa/y+e+2ZvxrJTHXjte1Ot7rlo1afZOUUxeIu2TMaKgyzAy8r5d5H0y4
Zzh48XLfquvuM4w0UFhee9HbKb8HO0SYNd8WCJFsVMKNe0vx8HIT+Nwj40wX/dEm9hCzXtOkewwV
CuJzvyucTc37mkaleB80QcFVeqQwdii/o/rsnTGzKfSiW4/A/kCM5XhvUpztm3iv+3CPCn0AOzJD
Q7WOjE5KWNas5HH32NQEEjfCAarvI2Z+x/R9NhqRfmnTMAJ5QbDDL79HsFg5yxwgTjhYGGmHAZGF
d4LsaAdc+LX0w+YK3NOW/66WyOAne9QHERbK7f7oXCePDyLL3C66tcHoXfddx/+fdTjQER3RhqcD
1rlOHiR5HhejYskODWPF8o5HLJpjf5k32bTlkvqjaDt04UtiqwagFX6HWOUd+d+fMJOqJnMYhfBp
9r234qfjdCcy0Fgvv0votflr1ochupN6N6ECJbjsjXAI/RmFdSMxqMe6d16S+79OI5zdBttTBZT2
kD9I7+xdJZN8LrCZiAQg59+gMG5zl1fJWzi2ixJ4VbhtSbya0kKDbXs7kMzVsCWdRjNElgfhDKe0
l105mA/9dLg82Os9Qmu5gFAuVIRc0yWpB4xveQaO70k+44/WtBwavhHPkmTHsF7sD9nBJJa7+dam
LwsLvB1gySkmJef7lSUP2TE4K8eknwjyiXHZjmU+FZvHzQB/IPLPHt5EFiIRu9iTNJKCaV9DrGb+
CamsjT2Zmz7QXD6ylnKcttu5pC1iQmbkucX7GiQqjHvUdzYWHDbu3UWCyaapuSwxiiZm2DODqQt3
Y2JucM7QVZ0rGkjJ7C/JNlMmmqIjUqEPJ+m5SCyyFc19J8ZCNOIUSnSeeK4TFrC9YJRM6wZhfL2C
OVASbnvdb9SsiTE/0WPx6R10pIbmwRhZ+cNdmKCGGNpLhlXRuLzFwdXPQFXhdSMZuZ5mGb7+76X+
jD9rSkNIMaga97BUgRrC+rijvuTyqhelOIxYPWT9iLqMEmxFu2YTNrHkK09XmbkKd7TJwgXpdnty
/5g345l7Gc7GnEmphaezGkwWjE2Vr8yNL7uuUTZIEIdeF3yyodUIUJJIT79KTu1YV4FY8/cA4x4F
k85RS22k7mEimcnHPyzu0Z2kwVb0Iupk/8nsJxbvJgRiGAtBJFa4cZKrNZN4fpO7nfonVzHlLd1C
a8NXzqCDJpyZeUzx9XtQmUsAXWxPLDm9EtjVXuWPxYuE3Z649/8ZlgPqy/RInmtUNBH/U/TzDV19
V72zYeNW4SghICn2TO6lRaz51XaWNKasHf+iCey1Fy5559o/WKXAj3LEJAdG7k3PYqhfJQDmSeht
i4Ib7bHSTstKdzsNQPf/RNTFOHR2WMaSPOQ14Bt5rnhqkWH9pqDK9m56RET1vQcqJrlqYxrf/laS
B1NWPMH206RVnlXG1g5AgtO+/t9Bq6aOyofhsUMUq/ovHKAIDsKwEONPafDKom+lEccQF0wA7rqJ
v7w0D5sn51QhnLm/WCuFSOLU57FSJfIWNBiAwpNQy5oiPUzzW4o540Ft5IU4iDbXr073CjXbyUVL
F5ZXUqIOtlwyRqM7kGxITgC9NryGCnCOBSFjbSeGbpMHQwNPT3ZJsV8HN5Cq8i0NNOHWhBD6NhLt
EADiqYG5jBraVWMWDQqgC2gm+y5aZ8KSuCRt6JrmdBzbTtjXMu1yYRyTTD/krzPNwXU56nkUCboW
xj/vGF7qyx5XdiaKPI+00smLkYy4B6AXERMZmE1XCoh2MayxHFVWPiCHs3qgk7c3DP/CEpBpuOZj
0oKDGD3O6obpnNd9S+QDO5v3p9cAmGHZXER4szAanTHwXyoeTR9VyAqE8/Ok7gjZE/OXTLA8VTDL
3i3FgASf+Fuk9Se84JbtRTzfDbiEQLL0rPKtGA+51sjCk73TsPQoN5VsZcC6QgGV7Vig1zxFiNR/
pI17VamJBiMKtUFX0dcwvRMZ/gU2zlydIRIxM1uyLpAyjvpV3fc5QczaQ/J3Ed12sRWzTcfgTTDx
ihsaN+okUugvc6Ukj55ic+DYGJCAKLkYvsTHhXZYqjEykM5wmQK2MeWP/u91c9u+/+yLDVWBBtRB
3daAx+P6F8hO+Kvb+xkDN7QkX+VcpkRSyLqhmJcf7BV3iHoY/ziJAizRiaYmA/ROs8mXfhoAo/MI
xFG4ljPZxov9anSAJMPQlckWM6Ecx5a5XrDruxWV9Nmduif5ZdXFXUV11EHG6WDGpc9974jXpzvz
cP4Hxis2HavuCcYqqwDG5zAg1yKVEvLolmHqZXCpS8bV4t16AxbtGECwExPPh3IXgAzhpj3TpGrR
zFGHGACf4NOyIpNKEXlcwrz3fB2X46gPx7+yXYdxgMqmXSXV/rWJj94PNH/VnGpaghZko8oRxpbO
OYKjcbTDdYKh4sBRrefEx+GcSV4iMEcNGQDO6zULulC8O1ycZomtBfNpR0HRSKSn7BR4DsusIjfm
xxJbLUErBt6wU7So9iz+N8sV6+CsR4iEmaiDrcB1eQfECvtAivbh+EZcolnUDfvNdNul2f7wk0n+
JjaKTMrgcUebZeXAoq2j2IND71hHdhdYyMuIKyVXtfXMn0lCEXqQdpz55f9RwR2PvGX7+61uwi6p
J0s49Zg3xWHkcp76d1co0Q0cHRZQKr9wAqADJCmEdpQkFaOr+x4AwhXuU2GPfo97EEt2HAbH/JnZ
Z74gaHxftoqSI9cc6e/p3r/pODU/kaGaP0pD21gqIr2vRzzs2oF6jdyJFTD8QSWmQrt6kmymVMwW
j/C1H/u480rX8qK4clr9k2XLxNONcaKEzwBV83b1GJ+ASjCqhsgFBkVfgi2Ij6GJlPDgQbjbUgLh
JAxwgmPFm8nE2bXkTeHPSL1z13Mw9waPGXHRoAOgukc9iQcjuLeM70NEzcp+aFvWBhk0hxF43z3I
oUSB1ghtANUzMqge1fPKY1+sTVvmbQjirahQPLbbG5HqC9YqxhWL2skBFiSxdJv53KdwcRRSD6T6
kRYB8Dmysg68QcXc6QkLwkQ3BuzCysuqb8XKPn4dG2x71THXEHm/lCRonqKOuQ4plAcYFo2kquH6
EFQkFY0Iv79Z855FyKp6vjJpn0zPPaoCCVDLduG4zlO4FN7FlPsJ/S/EqVcePMfWraEyt9aBQQyD
gq20Xh0UkOeNCXMG1zSzcr+6UZh6z1pJg9DLOHbQ/HUkZUnhfrg3Tb2yepRpNpTJwWI3K9fG9PLt
+uokB1FqB6/Eoo3L7eelBMxc7IQnWo1VmDT7s4xIziEHjXhjbjfvYscgZ8Fs1DgEys3jdzlr89i5
NcLSSicD8dbO/ewajr79W35oUrearHQpJmiJP+esao+CKkYBTIOC++zjL1K13boDZCuRfDt4A7H6
PL8yGXeMQ4fDBSWVftin2GarnugTWUMhb9gtOQ4s8SyBxeE8TZvk4Mu/vxpmxeK9DSynq/IVRnaz
LP5kvy+LFRQpdhwY9bqDfgT9Rb6p59Q3MdFWb+RVeDpYaSBpVRzz3fuNmtwL/5QqqiFuiTi6gTgk
36MtsveNLhB7ONkkmSS23avpLEukunsdF6o/7x8SzOPEz7bvO1uWQfG/FC39yTYbQ9dW7Zusi7Bc
gL7LGSUXTbJHPcr7fYk4P/3OjnqBTZntO6T72i/mKyvgZJ+qSvTKpg8yLi0O9J0uEwS1tgWq/+2a
g2aJZW37Ruf5kJmrnj0kIHKFpXTs6WRKS/BUJyPo+WeSoBKBbTLkmrlqGU2+R67f54ljHqYhiIq/
bTeupWlrzRQVy5WXNrYXFUu1NSzl7FZ/5yZbo9zwqXQn691yLC6bqjJ61y1x4u51kEmQnta7rOtU
c8ndA8tdgn+dUqzKpfJYZCAw3Eg2EAGVqd365JY6SScl85k2cr+WCEGNixVlNV+oD9nRyviCsIhh
ck8ldWNJP4spR2r2iAGHijJoITabOnNYTaZuzRG7tiqJCeNgQ4lOTLKBAraVWmY/MslWHDlTIRrt
4lFcUcvni3YgD7yqAdTqKjyvOhYqPsJEazyEHZ9KPxPPnI8WfTfgODdOuVQC0JCUGzvgRrbgdRhY
95Y8f2cRv51VrvblFtasHr3nnDHv69d3NI4OIPUsndEg5QGhQGJZizYDZDwOjTgbNq2ifCfg1Ik5
NQlPIRVHALucSrkR7b+iG3Is/foKBRvcrf6ftznPA2ziaoORcbd8mojS/BoZaWu+UyXlTaNaE8Na
GewdJimlb1FLchmjMjRmRBbqcyUO/7ux2zyQpydle5006KlzkDcUZ+Ak/IO+o/P+774IJzA7JYhj
qcGXl1QF4RUtw8NXufsefhNR66PZWZlUNKculs6V3Oym1vi6UF6BPfrR0wqIwLG5Hi+8iPB6YXNb
JelfjDA7vepv5DWMsmmi4mLDQN1ntvxOvQJL1Jt0ajjHFmGCDNKPtjIFMAN+xtJ+heN0MesuMI5F
9SxN+cDJoX1uU2al0+57+WhV/AwwFKoqZubR0hRzGwE/YHqec/wD971lzjVFCSc3mWwBlObKmY3C
w+tesoqYV5hXAOFbbOwpGoZXR5pDDPI8hf7DRYCzhnHa9VoSXimfiLIWAa/sYrPLxfHkeO2TCdGq
QE7rI1TM5NSsjSgLCfTlYvV77wmykfYofZcItQDDAxWkIF729x05YEc/NYtWchWOyPVVumBTF/mu
uZwIEW10j6ICLQzfPKRBLJCmRLDxj7wCgcR0jecTxU5jUQryguScZTCRvpXePjwVCXE7ptzE2cUj
qlJ9+hT6+oCE84uhiyhyIu1SXWP2D2oqqiTmtd7EiNWX+ovtol0IgoAuMJA5kggLHP4j0VCtdZOJ
HypyApTMapOt58Z/3DG4La4h2+oL5NSjmX6V6kJQuJWdUIALi+8xwAAzp6H+l2pwfXxpsRLEyEBQ
q2v+0HHM7M87XPTHnOTqq6qBh6e/WCPser8m2KhshEqhK96oc5kOuiVznPEEmQD4Dd1EI3sfVCjX
Qs190panmqBk3fynbZ7aK53K/fDT5QfXdW94vVLMyNMYxaxCWPLo5FWhDsv/ItbljaC/y/DNhi8B
rUF0GPr3fZVm+WpqfdnLKOWuSxICQ22RL932Fl3uZeTPWtVbNKPoS9dqcZ1ZhmpLc3jpyCOwWjhE
Oerpw9oIxw5vfchuB25x92zCqzddXdFB48dDX/xpXPZgpaOqLyn7RbJOpoxeLjOA5MeNF7sDsFEp
3rSiv1mTNexTGgecN47D/4XnU33C/V7U58DAOoNNiBXCJjaxaf09UdI9n7V5CuAeOXAX4BUbKan2
G8bT5mZlRs0vMUvtITa6KFfOnDB8qSNuj4rAMhY8EUs9gax956YeagBgotmZdZ3fVkH60va8RYDC
U4F/3Irj9Sr4Z/OZZqg2cHQ8X0VxV1oIvrsSrwVU6qAlysRFPxy1UKi9FHwZa69tLex4KalymEib
s0ivJCY9h1c6A5bsvl1YS9ZjllmveEuVqESm/m8zmZ3sYeF/Tq9ujG1uxEKgrDnvPxnWENPKxj2z
mUiitthpGB1Xm/0Bgyz2V3JC9O/HvuGj5mbEoZO3p1axJZ7aMQahs7mOLlEN4pUfT7w2JSo3X91z
H3L0agrVTp1dcefqNcMHzddsK2H3qj1AhUcWH+og8EDUj0/+N51p7HgreH3g+jOTNLDkYg4Oe9W+
3TbQLsvoaqmQpnflyoc62H3syG3AXvF4BMHJA8rV2bf7H3pYYOsj+tE7NNfjpQepRz0SN6woiaHL
Sx1a9dD7bcPyeHkCj2w+0oN8Mr1zWzobg/msYOVB9YRsL7YXHkIx4AQuKCOEn7J1FD6Xy5yTTT0j
GhBMVSwT/A/WCoQjDHI03EXf/+orQ9ceP88ImItxozJmTzxJ/Yx0axs6XQZDdzftM8/8xwG6k9JH
/Tm8RMQxqKzdp4Z0B0Ic6OJsJlO4eHfDoh/yyjRTRyqYuVUOTNM1JMq4ebrUsQPUtUjK4Vlf2QhO
Kz1If6Sa2MoPLR8K9ofiYbf7BznITqNftOV1mwhpT84pZ5l0tu2OC1ZPKlfoqagutsFjUpd9ACEX
ru57UK9XkJSCYEbE1uvvH+yU4m4ZBEozyck83ouSa0NG54x5eOCjpPBrt5HedTl8LzaQBGq1Yfw+
mjzwX/iuCE5py1OC0S+CSYeiM1cmYsIDrZAFhETv3hJTP2lSd7qsXVYel8gA9edhqcsYmgXFOgND
0LRHO7E762l55tjuF8QmiCpSIfevgVHIfYjpOFa1ljDmCu44IqUfpagwT5LCS+4u9HeYbFGDN4D1
qZzLjugMQp/GzHVxQ04PnvkMnv+F9AdtNDhZb+nQwicm+jX+9nusTRBBj+u/UlvQWcAAas3XT7jR
ow4jd744icVuf+lJf9YEclD7spA5OKLlMu6mWP6yQbt/9jeRSWuXl6iSY2B1HEFpMlgKoROzCH1D
RrcwBCsHb9ZRLd1gUe1LPnMdLGBw0mJPRGkYkLNYs/JBOak8i9aQcllmT70INhmV1ijPrWcoHyxy
QISagxRjiqluNU7LvNge0FIYBF4zM5w2Vcm0PlcmNQ1c+xDmOi6s34SHhg3oQxetG+aO+vSOjn3D
g87g6AZAr64uYIJOBTVcs6ahzbskx4rV/gQPlbrd9sammh2Clr7QxnHab3fHz1ezExFhftoc8vqS
sMmxQx+puWsdIHtrxZln2vQsbSOw41s/u/ql6A7F50qwa5SZY5Qux6affqQnudR1kctPEnNNJrL5
BrnGJgD7QJ6E+E0gG2c9r/YHOxeyDB2/YTo6Ru5lW6o/2j8ywmw2wqWiEz56MwCJbst6pa9iP2WD
HywOaVrmHrIqlQeQg5MIFSqg46DN68l3tIZvQwdS+mbpw2bMAGRWz4HYh5A1UGODRT7PH1pqZZi8
0Ks5tJ7rrI6xj3CkdYvwo0Zsge5U45FZy51sLUW4byw/4klNrzETePFdH9/a/htK6RpKi2UlPVKh
pHP3ZctNeYL3oq6+BbEXhfYq8f/8xB8VYXphtA6fyw6MM1m6Y2u7Q8Bd8JECyMKnu4x0m8NtG+mA
OBFTmh3LS6O+hy9vZvdUH6A+qqdSqJBmYwX2U0UQVDjMqGMvR3A+uVIi2+p+aRUdgwUIQzAnnBD1
qOmhAUf7y4LIL4JQi1TF7Wu13JMcew98/JRlC5VLeMhm4LSEtTTcys8L+0KknM/dItym+MvS2BvI
nS5Cj9CxG7cmNU3dMiyE7p63dqWRZMpdkmCfSIv0MMkm2EneWEtOicPjOv2tpCYUnB9jYN0X3RVW
qExrJiUGQx09ZPVbXoPykqnapAhbBr/WXyv8vtMSh2X1DrP3r+IdlTO1UGRFHp32ntkfb8Cg8CxW
+YWbFf36wGQQl4ftA6x4fDYBqfn3GYzFXB0FnA2TJnae2PmMJ3erg4+T/Le1Q1TV5Gvyhp8RLGOj
P83RAf3Yz1aTr8s6RuxIPInkXk/0aZlF6eyF0Ftjd4wzAdyiuVIaBpHenbeRcqQIN/NC3hiyJY+P
VXLpnWnIGtr+khfbdkz1oPiQNhrvb3J/J1VaG+PWszyVPFe1rRyC97ARqh9xYoYZstkFmby8wHSk
axpZQxqh2kOYPAIsB6mZr1WV/EnyBskoGugslgqojsDUYhbqu5UQNrTBjcXyR5VHo5A4TdMu91YZ
+4EBXLmmyo5qE0AHpPZ3hAlY4PdSqgU1E1nZeIiwnJURQmGjUeJb2QSZgW7HWrtscaKQrH4jlk3c
neHzFegviCm23AgA1xi90JT0ZJj3ES9RM28HneX3EJ2RscmIm5luqSjQwFxUMO85dqrGT+FK/KNT
YjhT/XC4/vvErx8PJcICs+fRuj1mJhcyDXMe1f6BXQHdW5mwfmf+D5i6v9xdccz83FqrIKg4hOAq
qyCcBmREChUHaky+bLiTJb3B5jk48bm0MPbWpugSLuXCyhAjIBkvpLlVL9xhH4T9jjPz3+3AhGTm
eImCYVZ7QYKeNkVIKwBuq1cZ+vxKGq9kdIRbaYz/ACWECHpFLgHMw1NpfKc5PK+YfAP/Lr01utL3
ACUm6j1lHJ+Vva0ohGjRUuwB5OBVob+sztjgXNVNUEOw2CP3bTNg2bbRkNd/IGxXAerJdVQUnMD/
IjCwCi570NAV6sea/7PcRNMjBKn1UKR3W9cwqkDND0If9ASNIo5vEt9SeYwxhA8B9Lrgi/tXQaZ2
TjV+avdNQmVkbyJ2LprQi9LR2LWiPVUgaVTe7wtQ202hu7MlFWrPltowvL58dYvaK5z6jpHuLh97
ChhEcfFkQX8mUnZzrbvLsCzdaL7Am8ufo6bXz69zSHHmPwHXVljKc6QdFd/i+a5VLBT2x8DtgTOl
5HMdbOcIx43nZGisqctMWJF8RWCFOoIQK/wiARh31Ql/SZLtQTDRyXGxlR0PR1zKG4cX9n5ygSum
j9faMC30pP+Ttpuo/TSNJRv8GWwSK+IciYXi4hpHhhqnz5RaS3/x6sFTgyMCPEGn1MN4phUGkPvd
grGlQaLWaucvCXzdZnflnOZa44LCqQGBBzic+j5SMTIdSzYPTtSwjpK0KTV60Ym1VTApqQM1Vhr6
yHh0p6CwzTnbO8P3vwCiMtgRxelwrupHXndpc8Soi72aCOa2q9knpSBw0nBmqhcqv/F7f/9axecP
NLCze554mQzncJvf6ltztrbPE1HkArURKtu7aBKU1vA+YZDxu/yDXPF7Z0rjYv8KDjtIJu9M+KmT
70Lyvn3XEGcHMCrZw3hximllZPaEVpuJUIDme7y3sxOSbjD3HRMorg2uhTjX0DRWsCCS2ipXbpXE
4sgkiXPgnokoD827NDTL7MxLuYwcby7IF1Hwhr6YKZlgz1QfRpNu+4lcEBdUFJ54jMhPvb8wpnKW
ukxWM7nAudn2GRSY94tDIXzYT8eMRPWiWGr9HJUQMYeyD60/mpHNp7ZrVSUTkVKg8cyX7dpUgF61
Bv99KS6tqbB2h36glK3ZhdPWHh67zFKi/jSIwj43SvLMqfye99cVpsatjl8OeY5kvk7iKbl5VJVB
dyeA3blnEMu60zGMu+XZgnNxngisoTkyfpXaKhHjI1vm6ybPw7z8D2o2qaCxbPS7pySTLkJfTL8L
qtvuGIWSwlaE1nzITeeHt2b5GwI2zUw89PKlAgQdEgb/jht8Xird/8lX2roJFrtEN9B19XxLrwiX
VPcz5zmP2OIPuBBW5Xq4ghCp6to0rthVzSkvrAkvxtZQh5Rx1nTizBOWnQIYbixbOC5WUTC5znrU
s4hbbsv6VLI7+jSGt4BbaERD8L3KSTC44yqKo619kBkq7vsR2YkIGhmGTjaInwjC5e/NpyiOFxZ1
G7Fhr2gDJkijO0G+CdYj7LVEA6oyz/yn6uZLE1HVgVyPtK0L/tiybdMaNJq3n7+TfQ55GF7ZVfOI
3WIc9uxApQBW7btn0Comf4ejXIvHPkUxY0DnGto97Q5UpLspTukQOqs6tV7233XvtA9q0rUarjp0
69Fk1DJqOpNTQBwrKF+eexNvkMpzahTo8rYQDOuoJ2239Zb17IBM8NnwLGA61ixx2rzrOpOA9Z3l
sOloHJt3p4VHKVF2gtu5ho1QOQy3Q/4cylRY6d3hdOvg3/gAfEEEWNPdt4Mufutmkw0oNAp4At95
TRi+VUOEzb6cawu/VV2YpJBxzZZ5IPOqVb6dRw3K65TkRCKt4krSxc3nbPzCjARANXkC0MA5yhZu
aoUOSfc1XUdH+ATNahQ+yDKJoncvHXvDp0n5NCxLV0hVgmIiA0NpTEJxa2FPVuW5Cv8aCTWaVM1t
JCG9zMb++3xcxStZAJv52zpRFXDi95YgWAZYDctJn5Pr+Ofv1Wtrb1elIBnfrM1cp8f42PU7HWIa
teO+8Wpuh4rQzkn0Eet//wvWw12POSu/jEmis/la1eKxXhafiqKvL2Dv4IrCR7sjt8n+eHuG3t06
F+/GyYniRh4ZrNWFP2V/4hLK1qx07xrSwc7VSMGq8NQWz2YPIkU5eEvhbLY22Yc/AL41jziiJZH1
JWGwcJFLCQSq4BYNsUFDdyAUsSKulYnrlnXEF4aX0tirNoWhtZP7dShSpuTjVYn+gWndT8PN2rUC
vaYZEZ8Kztj5wYxFxJ8xr1ZGcygX+taaFzdaCj5QD5PhPWJDwpcHPiHz3DiXFqpZ+GdJxepSqO2M
K6jH/INV68LpnOVCzJBNy/uF2fBMLPFVcPtosquHM3QXmxcdK54FtQ3/jGL19YOhDbnVbbJYVZPU
Z9PLhtV3xYAwPvFD6RTpZCbiCW3OF+LbTKO+TQAQIANNl5gBmKmFskgV4EKrKi5c2zvggG3qGL+x
v33Ik6SNdSxmq6N6sw8JBgRd6KyP6xORxuC75y681KmSi/7kotLWobE+aCVgx28sKvKV0jH6HrOm
I7sWKCbT88Xenoy/2XTI/7zpVXhFJQxCGeORffpqJxPQNTPf5s9gTx6Q8X0f/nZ7M82BgW4hIV55
4yh3rU7IiQl1JzYTeFl/uj/Tg/ifOaxQ/Q8+bs3WtR3o3YuuoQgELut56R57AF7cQ64MiURt8Ib+
AFPdZfwuPp+nu3fTGaVl9/WanG/b11S2xo0xgwjWkeQyMW5x8Jyhrlh91xDMfll2krwZm9YFc3gQ
n/39CrDJdXSkdJASyDwioFVXtwr4ujH9dT7/INGhMNaMVOXpfJEPk0f8F9LrqUlU3jUmhDGi3+zJ
MXMR3/y+N3ZTsr2w1gvSuA/7gfJTEH6syNnsnQD77qhNlgqvu3UKjdXDnBFmxw5eHA6fzPOXBfnH
7m9JWP2tUHVwdxf2R49L0wN9cAbDBgSBrUmzmZhy4dV3dllQj+U+6KTTrITzPX+dYJT82yglUGwO
MCvi8Dm8ND2fzjsZNp7FKfm2cdwl7rRgzbcs++jassacYdnrU+Zqtj0lI0aiSc2VD6Ew/WN191Jd
C/+V2FN1uow1J5RlU9pRtI+9eTLa3WKE61TKlpYCk6AIJvscOMyZhFzp+EME5i+oEMdPmgolvtg/
VABuyBF30iolfe4Yk6GfZa5MMrZlMu1M3q9w2Tg98lUWKhBRNHvg1lbde0jk5/Br/ZBiNT3ndVXc
KdYhO5aDKjrL4z9coymazNOubUsMwRHeofugsdriPo4tRPxTiXPbuJ2V8HJoJGjY4tvofaY9riI/
2Idh/LkwBW9LKv0uNDJIL/1ihROIJPjeeXt5P8+3dCsFrEEziKCR54KeU5yPmbB+LtIRvn/M4QxM
RumgryjzLH7ATJb7umHKmpwQ2tA4sK8uMVyroggrCGW2WlZNPeaxaf0izH7HrQRUTNjGE/K1LTyP
gZc51NIrMxPfUXrJt/CXXaLW8RbTxDO9hDOv+jvEzJR8EnbDa6cVpZ/3pgCbJPD1QeqVMs0U9Q1S
XWDqdROFC7sCol4xTmFErX5KaB0qdhwzRhOZpan+a5wAvnRMHSGbQText7zBV9KZ6+Nb5MnROdqr
W0W5HS/zsZdF022Jo/XEeHyFgAybsH4Hw9h1jecLDYzfFza4N0R+5H7VktJNjuMj4TCjxwjRwesB
ol5OMFq2SakaO1ZP8f9fL8Qsw6lq0tXSyDmcpo7yoOGB1k/odse+kX4lZm0kk0qQ6jNOhqEGpWFU
VQuej0cJLuOTBQZGlQMVksqrxy1a4mNRPKsO1XwsfvWA6h/of1R4Kk8pQ0fFqxWQmAR3OpUQrS0/
/XDIKJT9AMTNTLgkTibfUw9J9E6WHIN7jNHf3NXzU9Bcma6kwlkBW6q2tzD0qslOtBjZg5vbMcUi
/G10LSpSSMTKTjnhq8WydqdBbWAVu1WGWD5SorpimfyXz46UfRAvzqAo18/2C7pNCMd87Onyrypo
hl4fYQvXJmaVDuqRVn7LgQ5PV0vv8ZUS/wWJsKx6CC2cd2r/KXeM6YehaYPbDRQNl7Pp/a0rUvD6
O9k9RMAmeeXM2VcSS6ggmSq9ZCkWJ8O57sVsP+xhtpIpaefVp40zv7/hUOofG2f9w+7Jq7dhlfbz
uVjNXi7rUwfoXdFPTDPlQrz8qarKLVI/9YQg+mJ5OvXfv/qgx49x16AvWJ9DpUtOk4Hlp5qArqFS
UctjSjjzxpcOdAbUU25TVJvV9hvUD6YMHtXMM3BA4L88J9yLZ5bCECcCNqs+ZkN1xZ4a2XjWpKit
UMmKpQSr7cmd/IjigRdlqgi4jTJRW6OlPPga7R4PeaWHR05CmN16NGIuaF3yO8leQJaCKG7ZZYMW
zuBZqU+xSceAGoleMnjEJpgw4bQsDxpieNABWUHQPKaXknpWbHD2j9HEuTOIR+LTkIAc9ZvGEOXo
6XslVRxkWDWnxmBR26Y9LLa7DtSGg5otZUxw2fpAPJ240WW6UX3VuabI0GfS1CWcjo6dM0Q/6ygL
YxuZ0PI1JSFiPD30fXfYrJ71tqcgjMKJhzHZbFdvRRAyI1w1Laq/sFbrD6NqucZEAmB64NoV5SZ7
Vuv4zSZaGV+tSiuiGV2+nBgoWRM4QZ1JlQnRMYTk8Xom0af2Hw0vMMMtz/xTn3lr5Mrp0JfyvKTp
ZXLuEweZikixLw3AYJOP68KVSHfrgmsVbRxldRJfjWcXNivnO706FkOHVsI8wcKVEj0w9KHRUvVs
PksfaH+0FSfWoV3tGXNsGH0gcYfkfW+k4WlPc6c6xKOrGyCjK8b/uXsSZCKsgwiMf3TP54qrdBR4
LqC5/80bGBD4ripL5GWRhe9DY77yZoilhkkkHcdxRj91EsSGG9btxNa5/Xh25+TcKKzbt+Lqw1NA
pmEsrHXL8kvgri7RAbRhd/wOe21mYV4XYt36xpUyPzd6GQrbzIv9HsAjnzLtJ6dqXGJu5N4+y3M6
V5QeFL58AVkMjy8BK7qLRAXPYtfZrfZPISg6MPOM+ggk+B/mOZ4IXbj1MYU60K3RUC3maA1BCWjd
5WH0yx+KUMaXWCQpIcaBxd3SAlWWT52hkXjPLyiu4Uhz8SEVeHgPpbJVBSFpuiLtuBWFaGwaHUNP
S26DdSk/SuIH7wgcJSHxkV3+3F/0OzvTS26QfO7C3RSD+D/MwuxSUwN9iLLBXsl/jaqWo1u7vnfB
nexNgxn2LX76nLsuzbQFw0qYBBwmTTR6Y/tuTl7xHQBcyFItT5MIuiDiz76pV3wU0IlE01xfW+V6
OSz6L5GLLup2mCLlrS+/xcWJqzGKHyDZ5yghstFjLu6h1C/WI1wmjnC373+f898rcX/vrsAtvSxi
4CWVH1jhxCj+jzrs64Wiw/nj3/Dl+M2MJiAEMawACNo8SjgUInK6oJvypcf8fbnQgAwLSlTCWgHv
FvY5fkC9ryZtqpiaNHi0AbQxC39kVw5tAptPyXGMumLjjXfM6owBBQSUGiQsIcf/bS3m7AWFU1V7
WvrvJJGXE3PKvzA04jtCbD9Q0GGhHwQ8TVhLl+ffA+FvR5OD8x0uo4r3r8sNLoaJ3SIvkyGnp+TN
if79qEg+ae0R/dYr/9zFRl7ffCeD69Y/JsL3TEmLGs4P7VCQJ2E7qZE+dsHkFELeUPe7VgPv6YrF
8ETpcF7gUNbiSRVqiY74WtJ0FJ3scyXGtSthLz/XrH6aOv6XD+r/yOlJNQNEfmiIkkCXvDw1m55U
JdixIcFNUp0miy7F5scaHmh41Cz9jwB9d19gaoSYrenhygWPbJdiUJgYv/OBFE2qXmvH5GIMp2CQ
BwvkVrPe8RkJn+1GdF2juz4ObKtJ7I7AnQXmGYPcWNM0JlEokCvSDxw2qOItxMZ3a10Q6jEsWdYr
uQ2ezeLA4Psgq1a+/2Z/My510HHc8NoHfZV6hhw5ihPWEhNXuy9+DxOdi97azUCubIhJAHVcqztS
v2M+2y7NfkHyeli/v918rU//TwOF6kkWeziM/AxprqGMetUdNoCaa3LoLAViHfY/Ej+CNrqWVeBP
Mcg9QkESRfQIKSUytlZ7klLq9lte4kTz/dYpgL9OGMcNb8Bb9qaWd1qUxV3CdVNDwl4vsVvV3t7N
/+YYcySQ3pOBo7iuaRYfM10aDIia5IrwVBT9vE+dXJZLC9KtC3KHQAXmZ3m9TsYxKwA4aSMkQwga
X2iuOh4MoJ7/I+1QH0chdZJILLJAhGTQTD/SamPKyhOUDL9Fk2GXntotfk9lB8ihCNgJVS2nwtV6
N3Dp8AR8646DKLBNuIra/HSz+biROCHeK8iZ+IFUA1X7F2H/HcTTmY0gS1jjs68Oz4WuD9urXM0Y
NxrErk+nnWsX7yat9oKfS5jR+OmlxMys7iT0VekRs/aW0xRcmZwtq2zF1JMkmIC9Ili90wPwq7Ce
H74OFkF+NXvKWLi328hoqPjwy5E7BsA6avIJuhT2RZq6BEhjlCMKks76sILE4CcA6HOcoT4nn6hG
7+3mVG8Kpr2JMkm0mnsbamJQyzcdlqRh9BRLaBAVvs9ivNNiKwly7yL9QzmNP0BfSNA4Ik6orV62
t77m5eVuqcNUgUbuY4bd9eKkmDEy3uDb1+ws3X5lIpEn0ic31OyxTQZ7bpAD4EUDfXHsyZ+vKUIG
QxF7VQzE/5bBJ2MnVlHfJ2gTQ8QQMdCCqOJDiQSLdhKOWw/u7ih7t4779RwkaPakX2B+y0Cp/3Kl
+8WNjiAsG1nTqFbv/KORh9kmRd8IQV2pnHLvzIyPcOh707bjQDiClPzQNYB2mTpTwiZzPsAX4FsK
kmEhlhu1gbjPfe5IPH3C93IMB3HVlgmxvMpccKyMrv7JaaObCy4gXBXV3osF3Y1Lh9CokpXF2LrO
RQVsHn6UBE2qI2QjJ5ch1Vc7KaCrPvY7SSGfBTcbo4jHHV/NGENSHUe3SP4NHgAPfH8aLlopfSQN
8+KUv/YkWCPBDKRAIcxtjDoJ0C4glWnjJcgP0wDJ2GgFwVgE6fHjvvmcrxJ0xMghZWKscrpul92k
sUDzvykt6VASacFL8/FCTvrsgjpXtphow48TDZO9RKuK+NPNH7U0jPzK1bB+GbQCdB35v6WXAdKA
qQGajMABguY63yFT2LHpHBYIeuQJu52vcjBGgrTVCACNsVJ4WfJDp1ViG7mgk6LMwb8Iy1hYLx+n
LIZQzr4slVYgimwIfwEoew0Kwn28zHgOLGwnA7lbwNtO2JD4MdXrMy/+NGsWaE/sqbsad+oS+++L
v9DPVlaK9ejB6wh6894rA/YZZGqWaXYSLkovK7d0q0n+Paqm215utbDRNpwCgpuF6peJPms+zf8n
FxUmnAM5n7MBxTAyTdqk3JsmhvnbL8DTTYJA1t6qNmNMd3q8OH7cDPRwAEcKrbCQCVrvCKaTc2bR
dWg+leKfTZNMKJlQDNV169gGlUZ0v0R8/cvXMaxFC2lAJ04RpJt9K9WghhmsokKDzYusEq6Wuo4N
VXRLPdSGot6vW1PBv9aFblZkJ0DtyRH+3z7Fp33pNyHsQAEYFY+Qso8i3kuiBo03P0y1P3YslLNo
jH3ApbTWvmB1LNCdcDswWzT8hqNX7qOojEj8cQGkqGvbTiQUZgyNjAtqMQx5Qns0hxCuHdT0z7MZ
q04emTQ6LbSf3T9K6VfcKRQOAo6JXj+95zHtrSKH0VzJyB1LLoBFBtWujrSedLN8mEguzW/NBOu5
dogoarlT88pLjxbKo4uHyOv7nz+S63fAXH64O/r5ozmv6JXksruJlQPrwKTj71RmP4+NHP3ktFCs
BYb/RMDtXJ2DAXLNJB72YBFE0YB7zoF0yL6icadY2RALCi6qrZOBz2o524PSgENwE2lLg0jNcUnW
1C9xSpgTenQib0dH2xLB34Mjme5K1lhv37wZQC4TpLfgI2nJgPHFIjIfYgmY+zvoGf91g+SOkh3R
YHkYBH0ILFSFotwpvOPYSTYBsUQVmmI+uU5L5ErrA2WKnf80lVUhIQus3rt+bor7iso9YeA+HELR
wbtF8x2zM12gW8tVPdZ1x09/1PuPaKNxF/DpvbL538YSPhLrc2ojL1dVXobEEWd+IcbzY6oabIxd
AgTi6ovo/rlxg8Txzd5i1IXtDSNu24uo2sDj8GjA28p84urw6KFi3qqVj9p9EMTvjqydMlL6UlmI
g5Ho3FeM7KiCVuCA8LgfHIYXu1V8/NzayyHzIskKqAz1RlBWvU2rS4bSypBz9cLkLbH4TG0GRGBg
3sr2N+Nr8vu13lLemFnuQBGbZ++reIW+HNzR0aZVJgntC5xjm4sXoE3sRslKu8E/1rNKRc285jaX
GMzsRVv/G5vIfa1gq06NwVMKA8IHA/qisdFn9IohdpuB/2MSwtlRLlJNuG5xKY5FOemOMA2w63Xw
rINx2MO4TKEheN+oDx+g5lybyXaQGKxPj3KM55LEtH8i+3mnbuPvu/E8QzLS6rtQm4CL/3lzF+ku
ceCaLZbSA4dIA88DqEdHflX3kRs+ljGHya2nW9wpUyjXidY+xbR9/TQQfEiRxF+jm7lLUytxmZps
kgjrrqMv5CxuVeC7pGMeU3FwfDNm1QWBwclZ020a5imx3BzR4cyq4PDogxEUg1Ywn5eQsMg14J/g
sMFjHRZtSNOtfi8pjJZwLzvDdIgsrGG7b9/Irn//9j3tjzOGwSFOwOJBTtVlSZ5+1HrHyp7Hz/P3
tvklKIF9iKbHsz67iDKAhazptk/VgOFE1DbHw1dwxEmu0BNx1/jEYDHcQ+BVd+4AbN3HJLCLoQHg
GJCr0l55JbGLDX17gROu8lpSBYlGMsBJaUPZVexT5ta4vczW1yuemxNZlzogtYgrPzKxkCT914bW
Y2RN7x+ZM6mMUnBURkKNuO9dN90z9UFXxmT2loUkEO0DXQOhXC7HUID/6IrvMzfFxy2aW/SxxecI
RD+X+3qb9aYu6rjp74GjyHeIsGEhtRrJgf8Qw3k9fK6fWbmc3g+W4dpek6D6iedOafIJtwqpcarU
Vuh1a9CQfNEsIOLiar9txjnPPgSUZTdWNFGChaF+mYkaTt1dTcTYd0c6rPEjyN7OyRwajlkIbQ0D
aRR/J4MnKRJOmN3oHwKd56qqPPVNaW3E4SUSJGBEHKa3Kbe+Yug6+1dxYXcfTKdYP5CVweoQP8G+
iZ/zA/Br7UOgC1IplnPyce3ZDzdAwtJDeYjOZjMuA/IB52AZS4fUQNs+///ue7t8UIY1m92Xhz3b
XMpFNKIp6ciSah0Xhs3eEj1DI0JBJGxTE13/b/K0NtQkbghVQQhB//H3/x4A98gXdBc2PXcMtPcU
chQfiUZVLpn0xP2inArFt5NNy/ly+CmalfeWBPXvfNK7GHOLGWUm7NdFWXbQG7Nf7P5cS+jYyRxu
NGL8mHUSqRMfxvjr2w8xXeb9Rw2+vn5vPRBMuEMvm2k059emn4Oa8EWaRheCxwRi0zHCB7enYX8a
yz19kHSG85OngB8lx5DdLTTxm7ETTa7HEhl5xU1YqkjRrY0oXnp+5DLkwAW97DRCY4+AWBjrXSDB
VkTW0tzC+i/mSZL08VQsi7Y6cuuxco4kbd1RMY0dgR/uVo3pcT2yQAJMqJCpuyeWfdNM+/vi0fR3
TbReLfl5kxrjjr7zTNNzCVhmCNU2kcqaTw8ks0tmiLP6AT6swXQVtRkyT83LPFVb6BtgBonuZjH5
jjuXOJb1QZfdwtEL697p5gwddD/Q7twwtWwgX2fEToYiJ4TMZ7bRkH7jZ9VrdIskKkaaeEatfXx+
e1iA69joFuinZkSgqxXr+ChQmWdNVXkuV77Se/IfFMdSqL4Mdr8ySwVGO6kcdjZXusowamOm/+4O
Hq2L0wgrABKr1dqGQAhgn5YEJcaFvyHl6v+KHohexFux8f97ktXY0tPuyxt2NRY6PFhv2DzfBlno
xQK7aW93PUoNWEY7o1GssZfT+XGskg0Fw9j+qLVzl64Jd784aTVSiz1uUrIxzS7piYlabtMVUugb
DT7WAXqPWqWsDyZA7LyiKecOkpDRFBa3614jfBVKqFlTyGkTrq8aP52dJzRSgVJ4rKEoq8/RwQ/3
dvH547uklCxxFlzlbPfXN+zKudzo3v2PQjrXMETNjI0fr47hNXnKM2sB8XWjM67x1aNZhWAX42w+
VzwtUvA+KhjPCrjUiyg5kYmG1AtKFgPHKPzttUTY6Llq7rRXl1ImYvSew0hwJmYOjlZwG3JbQO3l
vRDMN5R35592mlNlTbYQJmgYLKQyrJsHZ1zEirJ/4IE0HeDJDPJJhuVbJzJuVHZWvm4ovOymVy66
OIxTVS3IvEUpbKl8kF4bP0HXwXpgIeMy0ttJMMLzUslsT5sWFXOBekHulovkZb8hK44NiNhcNcn3
45g2GIAStnTVYMG8eryk/Hn3dsmBaJSKB2C1iEa2IF/46k98vUjIm7X5/MPuEYLw0qN32OaSuUzt
lixikRdyna3PeGMI8rqFUHYYBATRzHmuqHTcDqiZUEg/pZvKYHzdJXktjmlel7ZVbxaZLcsijTYn
h5asQF5msFt+qwxkvLlUhYlf3F9eLTfhLGwLDYg8S118ga/yuEExTSWcmA1ZKipZiGZ1czR3DwRJ
ogrBA7wF2T2ZbcHic7KFEO750R8DsnvZ5foMisXjCnVdhlpX9EhmTr0laxbVcEoiiZLKZgzLry0+
tv9ROuZfPkaXVFqC+188uwaxoFDYU0sEdExLPBhfdz3AHlBp+rXNk2zOxAYXC+gOaOxnjw0Yr5uA
quSc9REGpdbRnjLHuF3gNF5Q3tbd4WU7raNOsnhjpKsO9cHXooCyYa2scycKmoR5vdaAvcUAMDNK
Um7jvcYE5nzzw+JUuA3QhKYuj2uG5zhceXMuCui9/BkeiUKRVhn7bnqPFtO2sQ/TRD+Tl3jdP15Y
Ht9gw6qAq9jVg/+TCUMeu7AyIzZNj/cApOnD42KCoQ1BSgvP6Sj8VJ33ffnAaqudXmEIgjGRNemP
8BVBZA+z4FLEt16J4mf1JuGFEgX893Z74R7pr9Wt5RAQhVj74DXuEtpVaiQco+hlN7xsdxzqpeZN
L3OfDdbBajSJ0sEKiUViX+nfGhEFzoRgahDZ8r1yAx02UY7AoKVnbiJy885FhAIQ5izxAvoxupzr
eFKokIA8DFYbfnpEmXXBe/kmBFWxBYfhEjS1Q0195RWlljYCDFN/sLMM8EGvVCd9b0084EhvesAo
6LniWhVYbCYmFUnTMvnyJr7rSrhxk2X/IoZ9hzF+NvyMr10H/MAvOe96khGtza+LDeAGgHGacK+7
RkU9VEyuLvc19oLsc5jqgJe5tYPhHeZZ+k2DLZ+GqHO+hAh8MKL+ji8MT83mbgUITyCoW/Hn4sBh
z8qjuwo+rRVJfDEgR2sZ1uMhfn6+2HeXoBYcAhJy/E+BB46dsmhnBeP276GoU+7v2Eb0teAmNhJX
DkK8S7u/eFfDBbTiMHfoQU462P0NHhfqk6iqC47va70s0ROxFSyVu6+FcAPKA0vvQXPpSww+uAR5
1O34KrBmBUqELwDdBjlFcjARGzzua0ALsYRB78A2FlvVF1ajTAh8xlN0haTNGk2hT3eLCIRrDK6V
3dwpmUeNptobHti0HdC9WvstSKTjkp27a4RLjtQRaPkQr0RcEoR6uL1z/HbNU2MNC7ZefPWujdOe
a8JBKWPJTcH3khm397bJbIvRolH1/JfyvJ/tMjZ9bkcBoQmy9e7+C78ubRZFpORgWzXgkaraMQk/
iQ9LK/k/6Gl8+qILk8KdYZShuR3umCkclcGd2nWs3TAp4AXJ97TnSLhAQuq5gyVLNffb0QhWDXmc
pzj1G3ITefDA8Uy1ip1N7g/i2xL4EqqTfS1V759ZVYl2sz9Xo263disNlTl+B/q9dA2ZezDCJJ3E
WQWTjSK5W+1t/FPuzqLlBrD1uY5ih0FeleYoMCYuW34TiUjr+mS10mMAO6J+j56VjzDh1hL2hFUJ
4SquFPO/hgvf8TkECAyqAf79w++IQ2TAcSqeXr/mcNzimkYsUbjn7QcuVU8GbCwaw/yjHDAvSkdH
N7LWLqZwfBOu81GgdBSgWIcXyAaMtBX12mKApTwMdq/9gPfDofqP2Z4dI25pDu5eE33mBbgwrr08
FLQV56cWc0sffouPhxHhLSw+OMMT/SGdftXfQQz7rzLb3mV3PMlKD6EWu61NJ/K38EnIRPdR001e
N6GeNfm3xA+nDJQV0sqH2Q4SF4F89zhQVLNJYtnvJj5wAx2iZHbde2eJTpsLrHbYHHTYPeebCt3+
wwTsEGVlfPabmXs+HcotLLDIQyWyfmc7lGOyyrZ4J1qkr3OjETIhpYOU2Lnxh1bAPIWDpJf4UFvq
uncvTdBxPmboK08KvqGjBMIVmHVzazCxGQKai76HACRQjOm3TASqZ9HgMER+5l4ktka9xNS2s+Ys
Rt75w8GMf00FUv32zoJTMg2t6CKu/ab8TijUc2j74QKZ30fHndF1LfzDUEajzLoysSRINMFXlx9y
DlLe+xspClxQqGO8cA2X/BZ3vs6K033+d2bkGIbB0rqg4V628GFh4c703bGiLtGkYlPo68D0b1Zw
EfwcMallTmPSkb04v+ki2qrmpmBjHa7rNOWD5PBbRT0OL9RPy1jzruJKfcxA98aXziM+ae7fCHnK
NMejHZjmPDxUdOKjEhun2B5DyUtU2wbIrGZrSSGooBdLDrY4slY7W7oF5jtq9ioxMG8tknweniZ8
p/SA78yN94SSD88z8aGcHkj05qZ9yHnxeOb8Ndemq/Ie5BI131xUwR+SBQFZpBHysfnbckHy1N6K
lRV5ExeU+lt9npqLd1BOlsVVF9NxYmUcjTwxUNmC+1e1ODys/bmhwYg4nVvJBmnhth01mccFaymE
YfW0DnnUXMr4KW4TbH6nYzgEFXqrqS/xhnCj6XhrpLGClIuae311u4zYM3inaSryDcvENzFJ1EEz
5eVwye+AJ/am8b8TKoiyXog4uXHUIjwn3voqbsSx8TgUV4VqGljuir6MXNpvWxZCuHJ9+R5/OzbD
bjxl8106XmC/8cBd6rjFL7lTcntFcUi4TCYzpkM7z7NzTuzivJBO8oxGNsPJp2oMPxlNcFVBboD9
rNBMbNudBIUyqmE08eipSqnmOyVDv9oAC5XmS0vJyWLtHdYlbACvyM5eYNzCJKmO682dPXn8wYVe
v9prxgu1doAIAi1VMF8ixcgKnip0zSgC8LN2Ip7jMcBeOHXi7t8YX04/PmDRS0IM7Pbat0S6LGIG
YljVQ8ZiPmMoEcuX+3K5XVN4Z1f6JUe5x6Pzh0yYj6ZrbqaWqfk9HhZD8tjIfrOqpQUJ4vybHk3Y
ep+KudxBkLD/NeYSZYboOSEEFbj+g4nmaQ/mSGfyXYzzvLinnC7Obr6ruO/ScHeuca3z4y1E3mXt
QYZp1Rlp9vzY2e0lqXCQw/nkjuylnVrew/f6qnHZMKxxH68Y5O+k7M/kmEC/qI4iN3CHNFqHpBtt
QIYm8FmibwmdKn5LOwKPgqF/bP8tNP9WaQAK6exuYKhx0nBPzsNo1TtsZYfaNvC5yfpP4A3KSmcQ
rHArKUhUs0phOX+gNIG4spYudzi2jqcxcTm1zW271Q7o3R+9OTdyZMTXtOq3LMH7Aq6V/yWuwS25
hyK8vJcyYs69kVRAmSXbn5pzpl/ldXdanMGpylu0Vo4Gu8ZpyGHbQuwt0HnRA86PV7Uza/3S1VEd
o/EEJyRtjS63bnuFaogCO+hzRJWz33Y/7t4cYniWko4JWnR/kLTjbjBFv59sCAcbXqc2pVUeMwyS
FYKSFlDIPbl3w9hMI3c/YH/sYTHQpr40FFiZ6pFxzuMtQ7XOEbJp0h/059qSBr8QoawenOSzHVzY
47TYAJPm+lxsYOzB0h8TVFQPrckZ8zeVtes1Qr6ybneJct0cql7xcdQOXle6VRQKj3hsm2LG9DVv
DGKGLQmTbcotWN7KKCVwE0gweD8aeR9U5KTXg7CWH5bLbwMK6/XYIc2IVqX0PoUaEDZxqiGXjmkR
fTDE8//DmDzQp6IiAt8dd16Qu7S8lK36z8y9mB95Tv+9j4SStEOHsfcOIskJgqppkdx81pKyIk1r
mt46ns0hPOQcRixSr9pT6AJdasG4Xi+M2VAzi3olbQocdgUevHBQLcvFUx1TiepbZAB8Ue6qmBHU
gr+6xsYs/dyeArYYAGTGw4PFwFXqD82wDTjRu5g+Ci4HQPKMApHxn6jLRX/TjVC7cMWrEcxupqzU
SWBF81uFrJl01qrZVLaBFJ1BhHanu06/u7N0VJKD8pTmW1ElRInqvgDChkP1uIAdhejyNW4jNYn3
iVvBAeCDu39RqZPVDPdzW96xTwkRS6phuRi56lFsxSrz4rjx/Rpd7uNFPCVRPEhJHmUZWv/wOIZz
2T7m3x+v0tx0bweAJfI28aI6eu1/nhzs5p6w3khx/hzDw1qdl21kz6jQjRwz+/bI/NwWEmSwj6Ct
HnstHT5S+nFUyedC4o7mrV4W4FwfUuWH+La8BVXi//sMhozQSOqGTMuwSiOampTeiRL032K8+NXC
Mmw5McXLD4SorGMHhPuYAT0at/xoJ0YoP4XgHfGHQRJo7m2/xt31tfQmgI00GzSXjVtp5b0uWMTe
uCaWUjw19rGvNe4Ul1J4iO7mOMWA/+uR1S2I1jLyRRqjk3Nf89M7xSJtSgplLsgmfS4WYWRd1q6O
+dRLlEQ7sRwZYxP4+AzlUm8HXkHOExuclsb9iojld7CoyoVlCmWurzrVm63QsZ5OgqCxnrk8mKHi
XZTqoCwp9DaoSdtz49/1SZwjkolrcLJvRoerfE6IvC4E42Eva0lRC681QXEhyhKu4FLg6mYwOU9v
+VKvxLyrQFVBy/fWdbmtQbfJ2DGNaOtcM9WuYVp6W5c/9To7SPcFbGb2C/43xrKz6LIQ0wmH7Yzd
itFhm6AKUQlUvsY3XiZRiRsIRepGf5mRLW4Zv8Jl+gYOYV/wOFKTkzPx/qVJWDi11TaZFNly9sLm
M4RSuZ08PYX8r5HWaB2aJybaHuWgDVgcIbNaOZyWyO7jEpio2247L+JhYLHqdBFoR9RDX6dItXTa
842ui+o25XW4u1JELy4f+5Kvjnhp7UGS6NIZdIMLYAktrLYRAWpxPsHgfiYhYjO7JzE8KOScKaZA
LWR92QZaVHmIlLngaZFD8qKbYsoPpWk92ubCAEOiS7mwp9x4ITv4khByCuCudFpc4RhUA8S9CIyR
+hshHh8k+d3DqHmYBATd/XemAlMRk1E85Z9wh9hPhAF1Qx34gpqhbI9G/POyfC0Bj78O2S6v6/OC
dl294GfaIhiWeeO0y7fXju4gt85IRzjPEttk4fj/wCUb/97B7YkGZB2QdVCAiSU+664wPgZk4IpX
eNAUxPQuwsb9KM9M6YyGb8jiWCexvcwraUnKU3cJxjns5uvr6P8XzaogbmRuSDntY0CoyfMbD1GD
+ArCttRS9I/o1136LpzBEgDHatVP1fNfFb6NEUOzTGq8GqswozVRSJzZvs8ZwdI6826uYWi/E91Q
bCzzlibCSf+0zU1RwZr2zTXW7NcqlFhuZAifwiawvlnna9bLA7SO4GnjQIzJX4N/4jBbZK28uGlT
6Xo95J5cyaBYGu0OFJ9/8P+smzusZ1I7eMML/MzDBCtEr5CghTp3NtB+alI/1ehAuSdyxHTgFnG+
iggjZZUmxMyHcEoD0ka/UCukEKD6L6uj4iG3T4CMuPKB/l41j10iJxEtdJ0QZGADxGQt9V9D+P34
5wgprEcS82fDl+7riz+F5KxhvauuHAp+2/IZJaHmxCbEIsb2zXkc+CgVuc6Y9ewE8Wb/sBcbNVXy
roqtK12iUtShmlRZwVp8VK9K8zk7sNlbovoVDKSs4uXCnce/4rDVcTT/MhnEPJeTXWUIdpSPJN2G
vyiGRm97Z7fOl25/AKeie7oC4CY3rMKhgzE1WZihS322tKP7W2lzqwcltTbGcxYDkeI4Z6RbS4+k
ajO0rS40Y7V2wU8lg5SHkAwweqqMpXbQX/CQHH70mTP41I5RcUGm0+DC1Q0sphdKo5/Hx2HJLmDC
2ew/R7SCECncB7GuIRv6fP57wgYQfTrd9WNdMW3wDbC8ziZlE7hW1xnrshF1lanTjFH4nHIiINap
N48FL7EnclzDObz1Z1UXOgCS/ePGAGi5nb3Y0rasWEmLKgdcjLJg3kjCuYvLbeSniqGHEI5Brqqp
6aGtILeYub3h4I2yfVdxT2zgKbl1068jCmvE4jLIn/+Q1UFYQ4SmHshhf2AC32OUr1oAzRw62FSC
qWOzRVTgQXncrUnYIaHgMGZNVWEm676QkJpss9VrVGIYQHCuBsfDU4LGYfcTANcJdozf6njCFfef
GNIojwkgMO3ItZW4rDPV/c6eGUnExY0PjQnS5kR2EoZryfVi7JmB7bupqVxEp2hyY7omUOYz+Rdn
CHbtkts3qo8tACxuFXCYCM/8h8wqVTUlGOFWUxpubNvIEovZ+jg1jIuRNpRFcLaVTyLe/o2V2znv
Dcw4Dz+CY3Y0EYB7Yi+EYZ1AH/AH154Q8eZSXY77F62QxFAPgjJu3NuSzT/Ft9EL+4I7LjGYPxbQ
HUKJWLprvn+UrqgXT3EbF8ipvdl9ljiH21p3bvKzxws34mfIOlbEvDEhSupRZiGYNTKOIPSRIzuu
7f+18dvvYvNn9q23UafvlExPlUo1l7i2Ov2ExY11gFhoRIlB9bypuKga/87zkF5oZ4Sq/l3lQyvA
gPTz4QAMtGIbd7l0D/vdRECU1aCBvCADZcYS5flKkDGBp+RWP0Z/0xVBoAPtVU8xK3/6lyA27bjT
muMsUt5m1b2/F78ghda5g5EPlqbMh48stKuKW77cpl/TMUo3TjCaaw09vuIKA7+z5uhTTRy9lreq
5xqS+K5aC5pMTHqnb9f/tji/7DWR7mZ4g+GVor7LDIeW63ZquSDxQtLtwPUSOvov2F0HypidRC5q
U5rg58h7x0L7Yx35qi7LpPVW+YnqImV/TWiHWPxawyB0jN2QzLPyOyLq4CEtxMCxoqcCAMM9v3o8
ccZ9//e1VNVc0Ih28X/o+kk076uXl+5Ej52ioBg46hKybhhcYLklBcudnuGHfBI2g+vdP3nPeUq1
H0X/nIe5oqs2VuGUFXEzveUPmbCTMz2BhX2rglybnMBOHCd0POIKkUY7VIzr9Ki6B4iGFY/dOw3W
oYoM6YXWpsOlwnox/YdTKr9Bia53ldpYRzeCt8NxBd8a5FNs76rsYnSNF2K6XykRvFd0SKlSYBcd
dVEFVC+u8N0ytTWtgKPSTqmgCwnK0XLhfByCkzKallEn5jwqjJaFtg4w5dV90pW8OEWJYYc9vtPx
TT/9Oy8V4N+rqgjJ+b8Gq5B92N20bXvJ4T5kpdphYnnkrTCXmi4qHxp19DJT0kqhULoCMbcttyvW
OEbrfu9i9r5mJZi4H150g8drfXdvu4DnfYHlj+931fc7NzJJSHzsC83YzwD+i/YMHQhRNjzlJY+K
7BKL2dlcFMULDwIJllqHjayaP6ta6cqti4+kPzhfK14sEfALvdxVhDfLQbXNWXhg8ruB3SEgdFDX
GmhddSMe+ocpKpiD9n6K+RQ9JbLEUbKmm8xeyjMmg++R+wC/3/e3+BHVzxEe4/cqv35RXIi8ZZq0
ZO6Pa+8WDrRw9aGheqZNgmtt/MdJDK8ifRKy6cXjrUWMFdJEMGAdirLOHa25eBpy4vGzQRxHXX0s
zUHQ63WXmNfXd2MepH2lPRLRXk0HYeEOuv7tl/+h4JirBdFbKyPBEtkaouHvQ2Trsd1aFMELDzRq
8DBGsMYCYkjwvubDDvzn8i0AImSsr1HgduFtLHRLwrYa+3Gxw2D6LlcruDpZFQ7XWjF57awp+vtN
SV3S1Vbnb65Y48YC0PuL073w1DdgcC/GSHFBy2GOzbRZ3r3lV0yeQvILDW/PGzPrZSZGnQhNq7lJ
UHXAzLOf9ohiPl5Cs5DKyJ/jwbLer49RSxCygCeJ/gnh/FR4tGCgrtMczAqxAigBv7nW1i1/r/7a
n2PyhQrPhnBcSt42uNYnmh2HYGDHUgaeCkjqxirKWs+txJJMS29UM26qBg3TA8ZDeTv3HX+6tIS8
xO/SmV2dS8kZg0iXDz9iIp7WufdYm8iMhOTCowJ07nliYJPJbNTrYwmLrIiPm7kraXG1Ln4ITRsx
7aGRroDNl9W2SCX4pqcxwTK8s3EmqBYoiHoSFHYh5nYfdztMIjU+8kI3Xe5Nb3jSR/O5qn3vbw5X
bbxA7/m6GWvDBmuEhwCvn4t6rthAQOyjIlJYkicwtyB40UNcV7lulFktvZmIqqwFhlInDkBxn0m0
LcqN0Iyy71iMgpW6dLuxLJbPaV545HuCIfKb6ZQjZNidJzuyjQ3GKiGa032b2tcM06HkvFnEORU5
MdqMOd4cI8PqXZKOb4rQSS6CERnWCVwHVURR3gs/SsxHgw1T+3uLEtE0mIr9mwTUj/xYYmBgMIvp
qPDrg8olnslMU3T3iOycCpAdtvaiGZAX6qXlIKyUD7afxk3692ltWmTX8wnnF1Duo9zfyvBdSS/g
yaPULBw91qpApvyautAeL0zQzj0t57KUyQND2S01QgYJrndN0P/Woqxz1hHS9BLE84k/FXk7HOzU
022nN07Jm1WzZPFAV89j+/Du0BGHwWc3SkeGYFAtVgwXvL+3jxRzlnNChmxbV579E+0SGlqayo9y
iLK+RdztCv6GvbDYafGTEZchuRNyu7dwI3+RLGhhZotfzUpeuqiSwbx5K8FFzzGWPxhhUFCXY7yH
HKN9J7ih0/6G4Waoc3cOS8V01WlksT08dxitKpLLtw6Te1krxEpf5w5xNV9MReXaqaido98xWTkD
jQ0JO3tsUOfRM3SY+YYYt3jHQvLDvUTNJ5/RETV5S1bNL19gcVJDN7Y4E5vMWdKsuHAzUexBifXe
EkSOGIayyGB7Sq01pli2sEzSIL40l6KLAfuTfr16yNvbTdatK7MLcNL3kX/KQXrq5HYiWveRu43D
X3dK97085xiO5HPnezQdTPLtEdBkwplnlKgEk4p69ITtmkInhZt8OJvDnnpkt0HqPo6Wfz/VccCc
FJr9dFFEgpRykRa+3NgghMbfk3M4en8xqKY73TkBjdnDXrx3xuCtptmXlkRmYm2Rly5lwicyvPbK
DQh22XpWD8Epj005xxzTk6p+LAyvmcC8mZPgZPQHiJkWXtgJpZ44/6togqZZR3qef0+BB5A4QC2N
BphPz5qD+DvXzNYmhLgIWZ7chrQMT/ozccXGQF4mPtXVTIEQVRtvg8l1BVjx+1EKF90a/bbpnhTq
/E6ZhfuABff/1A+eGQDheZa0/+hmzxiX1QQ01GbOlbQx5OV6v5vf61Md2g4uWre68tJ/M3t551W6
DNs+T27c3soLFzW0GkrQBQREyCg0l5ZycJYa2LIqeJOX14iZliQPfDiC6seT9LscKMjsrkN73/3g
SKaRBAI4yhDDQYBMZ2UoXIMa6Oa9C7+X8tZU+MA0ocCWp+lBRhAw4BtfloAYLPWOTCGdanOs6OsB
B0cZWKKOqcJdX67slux3+73Bgz9lVDsUO705ASGkueJKgng6vR4OeYUq5VqOKEIYA9/Yf/6PnFi1
l+Qccgqjted7PMn4WADKGVLYdva++bWyeVt6FIb7m8bnC3ohcI/WiEaJKygKlkMhuZoi1PGO6+2d
F2ANxU6YOhLFjxyHk05BgsOIKupPdn9o3rotVa9K1PA2WdvbGNkjgPsPMz/jDZ0ovVPsjx2J1g3p
Ckhdp/uUEr0vTa6HjmNqxVBt2uyGYnxq+Xs7xslUZdRRg8pCrqAzSpehVm5K2UjQDycKHKLN1Jz+
GPW82l+HDTwwB/uO+eFu4jiHz2Wt3P6qkyU3ZxL67iILwZTTuoP8T+PZvj1NgcBLUNqAZHqD1d16
Ft70FB42spkr6oqpJUtdBBQDlkPrH7uMfU0biGPmMVVddfRHSfFSQ+ZLFNF7StQdy3zDhjUK8lje
YiX+nQIN3888NjsIHwCWgKIeH0PYlqtjrnazGVzDra6npTQNLRjyOxg2i6zjd+AxPqYTJiHjwsnH
qmob/MgfTQec2akgrN0yxupZPspD21OyN7J5fp5xXP/H4ss3PEmDmO5Av4o/UFsPeUNDx+r9E22A
bB6zhP//RwIaEjIG3WNEa3MBeZ3TISnv3Ru7DKg7ocjbEmhV50PYICUUJlOC/2z5izr5ZbMQaJql
Z5CThBIJiaw3A9c3meuFn91hclb0yraZDZFZtDGK1rWurW9ddInvC/2+ew/JXxWkDuhLNzgPLxc7
xJWjbpEOsyeZiU8r2uaXY20p8iWoyGfM2R2DF7L0N9HbdGIXmKQxzUgmoGiMOZVOgjw9GHdw7ZxL
Qhi2MTHc4jzUGpw3I9ycjfBMJa2JmmxXOubxfw929Yd7hIa/ejg0qAYN4dB3jGef5DOoP9ZL/cqQ
5jHqyIk/hIEaMnPQEvEnct5UhrmJVuo+WlInak3lLf8qHXQlQW3kAoeMBXdCROtvcY3KXkTUQq1m
CaxStqZaJqZHuCtT+WE7d8xMdZ7HQOZI+V+qm7HT/VrObWbTI+ZL7/xMFH2Uk3N8V6WGwEKyiS8p
BpZUslx5yM41JMiZ6DSRMT8XkK+QJPU9DYeCiywccHwTqdWKcgFB0pqF9U+mFqVPIZf5B1d+tdrF
rU9c6DpmKeX1n2LAuXR+Dh1h6N1QxC02d8ia+geNwicR3XO9FFQs8hlzu1bnUPIHJ8e8eVBYr84j
xSnPDSyTwNk4EcSljfbQ+NfRVNuESRJYSLgd8UVEmRTVXv1qr0LdcDTGOl6viuLy5cqj9ReRczvo
3vpR+FysaXxBlE+k/xY3hOQiaGvumkzIXtZyK5ctv5K/+lM0Jn+VTqalgJ2KIjFieqxCUdhoWV50
I2smbY6iY+k3BkcKGaD+OJR2qYkQNzuiLiMkG+V0FOb7qJaNNzzBb6aRB/V/Fm726UUOwQhvluY6
j8N8t42oiXNP15ujWGooxRT+NbNzOdWPjLlTEcSs9XGSvxofZyPprCIAmuExc43QKuZ1bELNZJiD
hmjY1l8OfLrofuy0siT4iaqe0pD9fV3xYQDcN8IcDZ7+zxhh0EVr/dBL7xn2HkO9PPy7QH6LT7uB
OA2q28KhszDZFUdB4ntxQ9QrZlfeveeOJ0UaIkEXfa9quEu7bgcqhhySF7Xcs6WLIWucN9x66SBL
zax5uvgU5o0yhzJGKkJ6vLRUeTnJqzZwgwB8stfJkcLueou+dAMCVtJs94M94U6NPjts7WNU2LJy
7F5FJRUHZogXFCLjxAUOTdMznOLblqdRvebhNnfebScT/wxDg84sG9T+/aISNcgLAN6IeeZDejUq
in8GqWAzdq0OMJ1wPn4IlXN5Mae7ZP8xVClJGZqkLrMQpVPjbamxNDgM/LwcY+SDZ6AtCFM/efdq
Nsu59nk72GCrktQVqR4A2PV6dTZFWwGy15zX8XvJfK5pDBrsJILBMIGKpbDz/co7ge9Rq4NTNdFX
QocuwzsMI03N2rwh3qKi56zcPSkc06FUVWTeV0olva0FNRZOq0fT3DT9x3gcytF7egq1FsBqUsoD
LYvSs0fHPHOAvBI6bAnzITgFD5DlDdLU0BKwkAKvQSoFRIpUgkwKyX+SovG5dfLHqQvDRh+lPCz9
1a7LwADvpCD33N24h9wv6NYa/5fI+Jrj5jprCGD9bQlP3P2IxehoL5lrx7F8wNQTBefiV0H0XNDC
pxuuaigFptyxPXetxd3Fesgds40pqeJsBLtesisCvv5mmTVGKXNN2ERiM0ZtoaMbPLOWrRH16dAJ
pZe/M9rs+1tQNiIGotE9qmibhrD5AIUKvV8CXhhf8XMVZ/Of2F3BJeXh6U6JvW19r1C8TlJEagNc
9MPyBveMqhxluGVa3bLQfmKbGLsPoyLi43AE/2GnsoY0Ks9hdGl/OxORXs9dCmaw68jlHgel4JN8
LXbmjOzPpN9g1VrgMFHFBih1+aQcN6Ry4MtEWr8Rp/F4LRhL9D8zkaXdcBRkf3D0CUpiH4lIbSp5
uAohXWRDNJSxJUqNrYniw9N4+R/fbKADd2hASO+LSoq0wpOD5oi1LQ52vx16OiVzaLF2YhRPtRaN
ROJBeNrYnXvL1QPFzz5dL75BEo79OvYvXqEZJ38qypdQg7v4wYs2JApfpXork+nVkpHrdEVkV9r7
7buQNdf9Gkd5zqZ60pnWjkWq628Ioney7A/p2qIS7ItN/YRJhCd28WBvwu7hsYWEI2Pn2nS+kTU5
yL62ZQh0objWJPp2Y25DAwnCgnLHS0nTzmToz/im+Q1fmUyMx2xoD+ddDRxaOs5fx99TdQuIraVB
2dmpp01eJ9EQ8MX8eQkCEl/A/FQ2v159xCROuw/WSYc1pN+1K3mdBC5zeWiwYBGyw67O5+K63TiH
jadUCF/rD/ubHpyw05YTPSDvOCkFAmYwEhDUCqmNubse2akI2JceXDoPMYqhS+S8AWRGFcov48qX
tI99b3Q7m/NXR0IHlCvFPM+4k0ineFiLVBG7b/2RQtsZLaZgc3XnR3lT6YKgJHKQbI4Moqrt35fq
xVM721KkpkhZx2naDtx8TIy3FUuYMLqKUI00qlBmf1+xW5ap7UgIj0pa9bqaGeMITdU1Z/CeRPAb
PYiuD5dXI6twSsf34drlsnwsHXo3sKwZ+cFn1TVy1alG+BALdeAbNneBqwOxRQvOIDZHVkeJZ4Mg
1e2FayAhlyRuU7sJJFwiIVNaq/ueW2goIIu5z2KyhqdXv5f1PC/IUlCKUzk1tml6G86WP4qSlioV
kUWl8k8nnO1teMVbThsZm3hU+Hmnb6BRsDJoxd+fgxlmqNYw005wkbSejOzK8EGR9iAl0MKFFf70
FqHOa3bcq8D6pQ9xF7GtSebz8is5aUki5hXvS6LX650ejjlShAbrQdHm+rsan123Z2OZWO+fOO0E
1+idm0ELIylZxbq3TZ2vZhNIBOPXamf91AEaEbR8RcJp7BsGvQO0ybLi+NzXIKFUOG+Na5c3tVBy
sLG442bACXYwC4hNlZ58tk2NAWAcIqxGGb/A6okrD+6TrBjDBkVXc5QSCe9cE9/YvTGXVsjTPzB7
130BdVY7BSIjtd670RnXVr07RdT89p186i8r9VRS3YGKHLCmqBkJHMDq+/0EvYEYa832OCsFCv3u
pgrdxZSdWjH/s+zaP6a9dd6d8a8ZOtsq8+QExV/0dTYUMUy15ZXff4ysMXsdHD+mK+JocHOl6NeW
5QSC/rcR3dVK74n/lzBtkRCdX+UGFzZ82lCYLFokk1Prto9LuAWjnt4V3CCYU2sNQIiu5cmn8jmD
ttZOKyyq9kldyzgJ1Dp7evPcDiUb/ouE0EjGCoM5F8797lxCiJvnOBgEXGBArkhSBN3U3Gukuz7M
m8Db/j1bRDr5bXtietBS9QD1gaCtyIxzYEaVQJ39KZeSPw7B74HUovtOG3CMIqyzqDqX3lgKI17u
549BuqqGnc3berl7QIzIkSgc1CVj8ZG3vEkxq/9CoKgxt6hVTfRCS8LdApXYqhGfpWSJ5GB0v6eo
WND4tLIXSPFGAcCwjR34GYve7vqZ3AOFic07LPpfO1dYIN+3BS8fILcvbWg9mUI3xYKl6OOx5I4+
bY1oMIMnLwqLVOTWeV3dvzWRuZdUckOpL2SbT4ZeQT04k6IvQ/bFw2QmQCUtzXLAc6jQcA1eIrE9
3PDQwK/3yJaDhwSQsjEnsJs3h7eNLd/vtwknlDtNK+qrz0oMa5ERiH8jjaahmkdex7ROhwVAI5mp
HIohY2bYpRN84Wn4MpHdX1n3LGMhsXdADKaO39AadPOjv7XkbyMfkonjGxxT8sQUDsMXrPcCwCBg
l2pV9UEYohR0A6qI7YYWZSWID30Gu27UYKfYyqxybpWVK4P5gxBW36f1K+p4c9kKrr81s/KwgTS6
la3ZMROwlbFd7vm0SWWFCXRA78IEU9BtnLa36wBN3tWSBLFA9bN3O8xMOLPj0mvGMPwDfon+H0MN
fciFiwLxBYe4tLHuBQiyOii9LUzq6dTR0pppq3YVcizUt0J04lPzeZxVUKcEUnfp7kRG49aYpdOy
yhk8DcAIkZfsVsLOVtPP5WajtnGkN8bX1w231Ro6DmcsdM50ERfVrmCxIBK5PlaeHTv7Ls85YW3B
/RLtHlYxowljLTSZC+d5S1RV6vj4c9sBD7ORRrUV3g1OIETYfnnjceKxbs3zvWh0OjWz2C9XZZiP
hKjp9nv8mQ5FfDa8MqEsD8rHRNoBsXvohRM77btUEcbV1AY8jHnuo8dz5CYS8QmIPOcuruvJN1kZ
CqkS1Q7AHgqWtFjbe2NT8qEsd7+L6UrkNhIeMFr+EZfVup7/JfKN565IxAZcPg3lu5Bbq66whpCm
0rzqY3+Z7B5csJ8a3DzNpYDulkLZUpaNZlXLknt6zJwaKPg2NVqBGyfMD7qYwng/kdmkX4cQO7Jq
LHyCDfo4v0NVr7HGKQdKtulHXWgrLISM2HdunpGXKwDWArxthw2MflcPSXYg6FnF/h+MjwprQTZi
+//A/Ml2vvokPP+Xdl/ZqXMpPaQx8HXbPtOi2iKFX7ZKxVmXDaEXwC/MVGeAppM6RXGXTcVSB5dT
tKqmLXj8c7/Y+SQ++cKE1ZWOTW4OQdE2CRLXrfBdVakSlZu91bbG5Bp1VDrWpmFqZTM7aWke62h6
ubNklKKEXG52BzFYY6i/GC50h94LFU4rYxDRzEyTUCX4zgLHxgUg3ZnRx8NBJyMwNrHRAUr4aojY
RY1TM/dFecZ1MvpUyZZNE49T8XblkrKFXNntZntKOOulFyZCzzHMPJXcwmUUzn93u6L1qI9syMPG
sN6w/ySHy/rEG3bafpetYRYyHw7ATTAACnUrXLTse1sOIH7eb/THtIcz9upF93lGcypAxwalA8Zp
nz5gqjPi9589cknJq5wIu3zJq7+cEAZ0r1TXDW8qXk2L1ChVs5WE8e36QCH9Lu+yyNfl/NOK7zl9
5ieiHaIP815veZkuKx71znrAfPKePYQzGtYWyAZRTlCIpLWpXrRKe+sl7t4jGndz+R5n8BulL7mc
fM/BZHY+yudg5cUdzSvNCAeSqwNIXYoh3fgLq4p5HQNb0XXFEfEGgsmYWpQduhCoYFgRQtWANP3w
XiAu9UzthJiWECDFsZj1P5PL+iI91IunjzkQ17/ekpnYpZ1YlqUPTDnTXs5Wl3OLoPHS4PBduA6n
Z6Ym6DNKHVE2HRo6HbSZfgty/YwYmm6aH/5w+D9Lkit+f8Pr+afNOYo44ylPuaKCdW3aD9VsaIBj
Jh0QopyztetUoQM8dYkMMzPT5ItAMVKhGzTjqwMDqLzNiA+vQFljzIxKbGuZbipP6jRuSCil1zCt
EDnpQc2bmHHp2SDHxXD+ksdGyiu4Qw18EmFkSqegfN+Pu4rhHnK6l1on0JQ2kdMYSzoS/lRsHupA
tDTK/QPb40Nt9VMFCqWZkoB3GG0nKVDDNPjgxJQCgTsT/6zGMDcLX3lwFtt6zqqEZXSiKtNof6Mk
9dWM2l7k3vtVZYOBKnxnOekc9EAtdWbH0zguQP0YElv4ULcg1EB8IFuKqj5CVG4XKl727nkZJRdm
A9e3EDoJ+aAIjetL/Zlys9B+kiRyCgbsXNa0hMHTjgy+2n9LjEvCSZwXkU9ifa4D08WdM/H8HAJB
OmxpjIDHC0pZG5YFXaLnT8pKyMjH4bbN1GWkmGNOrwh+PQG/wueeObSY03++xe0V1a7Q1kbjHChi
x1RWU/iTSvUSKxLYhSYFJntQOzZt3hhE0u3sKbXIEa7NkfzuOH/j/q3w3ijqN1DH+NKDPETTYlmj
6h7U+tWmjm0IBMU8WmbB0vmZyEqztfkwf+Rz6FvYyR+FEexLNv4dRkGblUfV1x82xVWiJupCE6eL
aj7bP939bjb+bpPuAKnbu/Ch9JQC0mRcPUEgenffviER6Zr8d+qLc6TOiooysl/J+9riusMwhlTV
pAbmd5jkWNQ5qdCq1RXhV0ZuiFeXCeqIWJyYG6daIrBDxY2FsftZaL3HLMw+p+jPbdkls6UGM4ti
YXK02Tz1ivjFBBGOXlfIua1tAfc5joX21vHGaE9jtF68S8zh7ltWj6rwKLT5/+2tjOOZMrMFdovv
T1Sh9nACr5xSovCKLn7Js7RP748lhkTOpqtVyzWiHcphrxxehOAnhjSnbdZbzBci23U7cjs5PUCY
F2ge9Puhu4lVhL4zTYYxLgxvSwwt4dC7SeUqBhJv9vppnO/1NRLHSobhTRov+vj9YnLY+/ERivPf
sWuRcbDHv+VrdCou1mFR5N/F+YUxPxQMGUsNF0mJGt1ny5NGzjUCWEVScdoon2w7PX136hiW57o9
ogqsy30QE+7n+vsExx1zv9KXccxQmeWBBNUz/qR5QZlfK3mvavc+79lWSma1SkA09cV7J6P+MUuz
N5VpgoX5RRlFRVP3lG2ZvZE4w6LYFRJVwNp3feK5RbVb9miF24HRILrX5MTPmFsb5uVA45mJpZds
HhG/eWGRZZsS3SMHMzvzte5+Vj5ldQrfbS6SgROcaXlMOnKd14qgSeFuk7DuJpn+hbCAkgTuuuZM
cAHvntxbJ2VAoP3ADwzkI/lbl16n5g7wBGmtPGaYwC65ZYXqzqO7N3s+/2+G03FfkzUrzgUz2/l2
eGx6E7jqAUvrYDX6+zQ6yKbiesTzLMMbCdRAPnVDHWuKDe4OBsNcQzj5rN9pMrm4d6zDRL4W/wiC
iY4YPK6WCQCin4d4SH/fwusmS7TH/khHhgyiTyyyQl/OFVbL0DqNOwqCRt6T1++6canqx4kIF+0o
SIowLD7yv2IHfNvyElFcm8uK2obf4ZFyezu4SNM/uxgyYqige0Z9sjgwCWnDbxij93DAgVcyWhye
OSxnWSMoHKzbpPsMrop+zQss6Cge5I9nsDVlIdEQMtmRN5vBQTlP4P9OriJASr7BEAp5Gfiy0oWG
jffP8tbrML0ITsa3r60e+wiPFmmPM0zkv2j8zxTQDsWwFqx5KhEp8V7spMZBBsfz2sN9DXnzREyN
buwvBgYMtlvx67a89SPreXg9KlqIfeVIo2Bcq01lpDcEXUMdjG5urs9WugJxcMden2f+gH7Q6XGg
XST2tP6I165mfE4tzvTwKsJEdl06JPim/foUK+Bv302wv3sWg3gtNOaGLOUR/NTRb7g5xtvr9k8w
LjjR5NW+H7r6D/ziJ43UAHTSYq0aUhwLzRXHqG5P2mgQK4Km46VGT/V3twaspiq4KaFfXl8ql9a0
gPmMqt9rEcpgGvttS4H98NZWQNvccJVXYiJojvizt5GPwMFCwByM2NO1Tx/q9BrBcqbxnnUQ7CXB
ca9YOx7SR7e+Js+R+xdrkt6X24CJzdj5svxARMwD8qdqzVR5BbZvlUhnySrEvZCUAQOjY07Zzvr1
3+LNnXllOaJUALmT5m87ulNpUorpNmKfFRUW/N0TJlr6+lBcp+JbBgkyDGsdICdC2lm65cLw5reg
053BteXCh9So74sJsA0YVFA5ZdrZlKww1E37+rcBGkP69v8XILKhegctkcqD9GnDokee6jfR0Q2V
ZNZ2ZdkvQzyknCoDeUOQc0SdwMvYQshS05W3qNV5/2H7pDLFFU1/oGoTev84KJXmwk4OUi7SvvkZ
47d+k26cS205venN3aFQrHPVqpFO3JL3TAbmX7VlheS32E/o8u+ONANSYgZqKNXwai0OLq3Blpm/
LdpUj2a3W6ifq01719Nhl4jAOJVsKbuy3uTf3EdPQuu7fY2AghSokVdDSL05fRUvfUJT8/u+g8jI
9VDGFX8wtDJnsbTowOBI1VWQ6OH+XMrX9aJXaExhESZK4XHS8WC77Abuk+8SM7vuIpi/9pll72aE
Nz/gab7snw8tfFLr4gfWxZElY0ta3LaD1YXJu+Ni/0IvlpiTl+lfEqLRoNqy9WPbmGA5myMPQasI
1Y8qP32PbYiXv84BoyDj9FytO/LTIYRC+vpkrVmOmtDtteEKhLHiTl3F7RXUBc/mez456vIbirIM
gLCtFUDq1TTNJdRolq2RBFr/VNxy85n5DHVXq7Cp5KH1OdJMCX66hzbJHydpnR7poeGTTLxFPL90
6zYN5uMaTZzM1csMej6582ODR2cFs0Snw3w0xd3XLFr+7nVzG2MWgpaRN0LxGC0UD+KZ0YY22/n8
vKq21ONagI9tzeEOmf4/H2MDq/XE7U8weCXtgccGImccbZ06xhfpq97NiE1N3NrjztenmW/KYvUm
68NdDnyP7td541FCcDUTRck+lmhrrNUsSjAXh3eU2fnw/tYcFi4Y4+K2H5v8CzxU/5ZHTKDeAxl7
Y/dwcCzDSNMTR9uMUt0LEAhxhH8smjZ0ReU6K+Gt77zKfswlcH4PbwCNxkEKonMU7c8rjTsSREL5
jdm6VJVCOtTAjCjSYLD3oHfYIKceANkNGTTQm1xv9VhP0zNBC4fG6LCFWX1dOxXkyXgBZDYbmzwD
rJ5T4x0hEqHk6pQY1lBN8TntNhHCDJGxDU+ZPsng7gyvMs0AUBjwOCmtDxcHGlcaZpmRihmuEpt1
ZclR5X/qfTgxymwCwQLyVpTH4lGY35Tl1yqt3Zpw+DD0RGvPosDlXXQuDhHocMGdxGEPJ5D029c4
xSYqzrviDC8U/kGSmX5LIKimf0nYHIZ5KIRgz1SIfpkVHEAlXPgSZQPmQV5oqc3WFtV5SYFR2jk9
R0kL0vXrFTa8cojRDaHuIBcBBsEqyv1lM6FlH5BkhHVbRsO3IfafESBl9RvPYAl7DwVaQT5QUY/Z
ubPymSIysgfd4SB9C7yaL6/+U0XSslJ9LeVRtrupv/sljoGOWQXbpUTJCspNtEeDxTS9G5vpm4ar
wvmrCOIK2sZT7jdFW0NChrWj4voWdadCqrJ9Ra6fElyZwDM8klZfTr1Zc2gWcHaf8R29w+Hc9313
AlpqlAmlhGEiE+yCaEMS13Jl4BSrPWcNqecjiDO2zzig/khpzuqzhY8UwpAYK98yfyw5DZJUQIX1
s92iVdt20KTGXCeThCETGgqy3hGQXqNVxj4D4V7d2tSFCoGJ9X9reQDrlVRJAi5v44p16LywYYMN
8oP1y1d+gtVVSA90JYt3PJb8yOjAxUe9PZMPMSq9/uNfCWjICFYQRptY+mi62bJL6CPvKiozv06/
SoS/aYUoacdoiyLojBWkVYfB3u9rlKCafX01Hjb48lcxIFcNKLM2Jm28O1yU6TitxRpIVxtXJO5L
pVEREPniR/08Ap7IcsWW3PnOudKmnWmMZAQZwyZVOhTI1n8uw4mLuYE3RgtPN1Zno/6dRGjXRdLN
AbwywTtvvpbzT439jGuQBJVHyF0x1oAVZZgTgP9L0teeyE07AafdcQeQ2mWjVGmy/rU0uO6ExmRl
zAxYrkgIgiOXDwWDoeQgXlhstJpRF0KSNoDR3G+LiGo72BXZ2mHd+9IiGVymp3XJYD3NSkgy1eMz
xXyKmev+/sXHaww8AcBJYjr4RQ+XJBUqqU9TfK1wqg66El/zKLio+MG8EaNAcuuJGvXKFV2OxSOT
hrAVUP9BFyXUovr4r2DCYfbBG+P9NCiuKl+Xk864aADBHxZRKcpcMJwFJYvwxPyvFeZwGyPsOttV
YAILO70Kuw5J5KTwwza8cU9f2tj6DWXGgN/RB3Ok6TnH6G4xxxZy5xVsp7oSqpzTc0bBntTy4Chs
qFlUU0Jcy7lv996WXXc8quX9s/Bq8SPdorpqzov8KBsuQ0zuETnjth4FxoCbQIih5PTmJCUciYmg
uv/vykxulg0paqV9XZnchipfbb0eGmkoDAqfoAqey5ANhQnM/gmuz3p1vk0+EXVKNnEYxKfBqjC+
Kv8NKh/IOUoX3QpTkDlTOPCXa7+7eUhvvTuvJ7RXuOmQLBqnI6AvZdaBhBjGxXKgyHqYSf7R26GQ
mN3TSliRX7ZL2A0ZCytIM6KEwIOFF9kZBOUbyXjJlaKzGAwuNtt1awGn/0U63OTbiVcxk4c58sNS
X60NGMTQ3dUfX2+UrgWFOazS3CkveEcsHDOkc0QxeB3rF9PBtZeszYAwoH8NBOOExz9DcIrgL0xP
AGZh3SOGW5x/M7W9ColHl6q4WiI1bUe7eHR9q61Hw88pYCdScR4LCfjxH55b3BcDdMjVNFiVh6mO
4LJcNAoIMM5gCEYW1BduMdxecW2Smx918gpo0lsPM6RQCxEfIwoAO22xw78HfxUq58FtRjTWV5yl
MCBxpMlUyJNhMJaKHtzgH0th/pToTu+fBVFfAg24vgjbUtVsbYcECzCoftg9AEUQXhXZwwqmXXlT
Do60u5niiiHmKyGwdgitKV/86YojtsOt8KJZUmAnLEquXatqQkri+eWJk4jXNiJMGXprk2OhYI4/
sVw/geR7wH4hmZ+hL57XZ61lmnYCzOj10vN5Zas86ekOsRpteqwqk5sOJ27xjgHtthLN9/TiD0m7
dIun1e/Sus2MFk1sUgDZ+BBEPAedaNXzGT90w8qBad/JDuZuyPVrkOJydoviELkSAzGav52ij5tr
Lnjnw2NRGvQ5tnrRb2A1B9JV1Fi7bWjdNDGomoYYUi6HhoWkPAUCAFyiL2C+yDQABiK9NT1P1cuy
hje0XQu8HPuk+Xgcbq4S+1AcYfqOEwXIypyoKECA6VRnUNKUD1XIWSpKTdMQPWyixVDhd6QVwPGl
JluGaqlOpm9nXXfYBs5EvIFA5K2y01SFj/qvGz0HBB1IDV5vU5ObBgcedh9fOzfe6oA3W0M/FwFw
JmzP93vtrQrkL4CjujB278JI+o49D/B/VQHWb8IdBAqDOJLt0XFc2lDN6x8FA045nBMtMHbhMSO0
m5EWHgjZaHRTGW/ngDLG62NhXstbxqE5U7SXUgMGE9SdG6zGiQGy6EU7JM9knrkw+Rqxjgo8JRfW
+dfLUtU1Gu37YOrhjp7PlPsV7X7puvCidws2Q+OATM2KH+UUGGWNsoQFiI1bqGgKpg05ejB1p30n
/ReB/2O2eOTh1Eilncri+51t2COiMAQjuOc748Siv5OE9wdJvfa/iBNBb6dVXcb22ogRiHK+GiUP
syqPD7pdL3Im/epWeHJcr8/amxd99HIETaISoEiczhZnTZQW5DEVEl4whm+KWtG2bCcTsd77UPAH
GIJtnaHnqmqrGMVseEF8mPVYgoKu0NoI8XSNnAydE5+rnaafSAGmUCqdszmZGl6h5bAg0LGwYCJa
A91ec/ucyjR+xjB9RbTeeQfmWif309uTY3gK/jQmrGcfoudkTpEoqrmxPlskOdn5OcJhYWZxqjnx
De39NJjVQghblF8tXzWQZMe+RbJKgcgfjSQY7q/y+ZEo9Beh9QtWv+nLDSBBnr8nwj3RfyzkSxho
2tBUvXERpjidAE1SOHbjxPpaXfEWKwI4Jn2ITYdWio1ZieM7PQ3UPf18amy2jXz1XrQxffncExd5
IEWyLPHZebiQtAYGaj1+58khmznKEJ8m1DvkAJk2goH4sJ4KIz6SZgSqmuaBDuoTUJ6TVpXCG42z
z+69hpEB7rv/17CEQtF+p3tj6xoC7rvfpj6jBpHDyp07CdPy/NygF7ieHutTCGuQWaubtknskMTF
0i7hzlG22r8xyajHH+xQQSFjr2YZIWjEdHY5HlB6yufeOlNj3tQzdl0IOKuGzSwNl+9BmgF383GH
VarALNlA59J5M35pMUSJP7jaEe4Z/c0l5bUSKXSEOkaWxbe55F8YRKCoSdGPusTCl4VZxyM9+EXj
wYtkRi1FjVP1ew2JB5hJg0tTiKq1TmVTgWR+Kx0loI3ez8y6jjCiNIS5LFOTR7CrvLxKKMTrvJPu
eLVfYffMRgnP7LbuG3wGv8MuMLLqddtk689m38A6nAboKJb0JWcpYtg0MV2DlWjyntrNTd8FP7OY
7WRlr2++rKe9B+/5B45Kg5iMe/L3L2nhmo9zlgU6O/4OtuGOqGVi5T8ibjM90yVPMbfM4wiBdM4k
AWqpz35BX7B8/cpVZgLlNIRPs4hSCKlPAZSRdyvSMTBac7yykaBIGP7PM55mxZMbhTQCPCwmTkbZ
RnggwbHX5uMVxXPxqydPja3lOKPLtWvpjWsTwaNPaheW/cul49hHffwDFmR/7+A3R1IpljPd/n9l
rDTrb1uZfV2rKgtSb4YmxuBDPc8cjezje/Y35C4pmDwamkXc9lZ0KD2lU1k9e1b2YcD0uAhVFi2X
8GTFOwSyrCZz6kRxOgMPabbNljAfMwpa/pMaqNO8wRpd0gKG+Hbv3m9uuboK8CSIz1P6YyYs+ICA
a+2+nXnIRkk197uS/9oYcWvaaf2HJgbV0wcJP4NnWD4HvbTLX3FORx9cuUaZaKxMkA6E5J6nnHna
/RBce26aypXd4ks1RnxfqTVkSGajttNHiVq/GKh8c830XWCgK20Vpz2IP2u0aNn0UheW10lZR59/
nsGPBg5JPMGcYyxHnL/21P/9L1SQDfHJTAlMNjXVZ8RYEQmXm4AQ0jdrJT/1jli+aAZkKc8zX2qP
0YF8v9S8QOLNSiN6Jc+fOd204pyJdc4fr/1LO4ddtH84RNWYdDzRnPSzG53+ZWIUdUq4/opy1iVN
hncj9UxUauH7mHZZOEecGlAWZoVWlgUJ32y08LmnA/LpJDzBmG2Cu5XiIb0FArJGvyeyowqqdG8H
uqfwC3kLpccs84In9QoaOhLfUqKRDU2UQW9FGZrFc4CfSoOSBULgrokyWKKLdIOKh373xL4Yxu5i
V58ZB+kujTjKjcu93IFdpASca5hZMyRQpymX8SkjWUMSlNbsXVa3mVBkp0dQGZaHc0TTpf38LeBo
5Plyy/Pc5J6fVewYYME3fUg4XKNPzYASDxKxxum10Z1UMH51VeiiDvoRQNCMm7qm504bYSOFME4J
C2szPIBVVHq+Iq1ag+cJnQz+A9WFVIZ/sTmu0hKF/6rgq1UB8s71Ks6xiC0MoMaUxg/V+iJtZqYK
WsHm8SF2/Acbwzjm54PeggWfrqdnq8BQg4M7O/hebbm/Gj++gXUvUZpCZCH8/eAnOV9B7d5C+CyR
3txF+ySFpMuVW8qy9reI/keebZQSiXTe5xUdKHDCCXTWWf1eErq+1Q9kruvvDDf38am9NVR4XIbA
ndSoYILEp46ynJe8hOlB5dRVl+2+tNG/uG6A7AsPx+zD9IObHzhzcnVJM7c4PlGcC+DElJOE4PQA
CzusePqaQL26FQ8D+wVleYwEcAlGqvDdxqN3X4icREXWusiknt9M3hG1KBYEczNa6KILtRTfNmf4
lbAHF+7PpZ/LZf2K2RLeNrqgPpI6cIEG+plwxqlX/reNWBOmVfVgu65zGiQvAs26Ffrd4jSIEj6z
JYxVtFR8osatDduktPCZT4Asu8mnpa50JsdWaj3IL0AmR9MSMd5G7hjrxkMSAO3Ov/hFPOhtVp3J
6mBfSe9nPswzMkVMHmYZ3NZ1VnQefm2oeIl7cV8rAqsgoftTkGQGQFrmaNkJ3rcDVWxcBlU4J6vN
BPcLBpjCbV4JgP0RW8YavPSLGPDw8LXuYnrgB+JfcVTOjdsxdOhpjsWmlkdbLi+7veAGvd2edxpj
OQCGQrmlrllosNNAZPq0XJ99O6jDN8ZB6u0KTOgIdpVzFqJjLxxv/ItGwP2o+TJFbuEBBAIJ/gDo
CuIf/1XL0V/Lq8txmRMpArEZeAdPDrdHBoGoBsFGY9sjUR4FtG/uXiUPzFmPKZqOFxcctmHUzjw9
bv4ZUcDhzgRyAAWBBMqteE4en94p42MyMSltoC/uRidSuov1I8jDU9jDO5KHyGS6egulLUxPug04
QzIpQ7RqlLKruSYGIkUx8P/WKx2hskrYvPSG4c2TarQNDfnlH7v52H03ObC3fkvAh13YmWGF9sKZ
taEfvxA26bFBX1VxKTY86Ls+rhHH3yvkmYUtpGR+962iajDnkwzddeCdeqEujB7kjEx9U3nvG8W7
jJIXYq6MJ6yrwCP2IsbqhLixeMXzBsfgiJI7SSdEAEpqy72wPc0gE44GzVo1v7uEhaM56yA/N1Rw
SbcyGgL0xHbJTzQVHpy6dNIU3zTlP/ojuSh+296TmAdY2oB4ah/SPXf/21OpnLv+b0LqMGjq+7EZ
dfT150flNn5UKNFn2gQhnxVf8ULPRVevsgEFwDIrxefrrjj2eQPyBi7QtzvkZmjb6pB7uxYtQ1Yq
gJPsk34PZ1Qi+UGxxZuE32dRpL5r2NUpemEj6Ur4UkteAbmeUzI4Ay0KOrSmvU6gBHK8IrOilJg8
QNteWTdNSYDXcNfu5dA7T3trmQqsTg53BC5MfKa9GdA/rGa/Qed+YHdOulhlqIkMsheZNWI3D0SC
2Uqqx54B3IKCWs730plGDVe1FHHvgXTrqWTzSpjdI2S7IsfFPQSwQ+dQY4P6jXG71zoUk9HI+7Sq
RfLhv2HS4B4jFg3j1LXRxb2WvEJz5IdXQ66ySIbpjQp1b+HknxIn1cMEWqhNG9EgBlZS1GbB5YRe
CRQU/q9GyZ0gdGPbhwH4rl+qV4h6haQef+HtBjkrwVLLutFv/h/JB9TVCAY9xq4Fl6wuA1euSXhL
hnxrwuIuhost9dWnsLU6pOXcOaGUXsXnHavrb/Ue9+KQFHcZe0rbIUkUqY5agf/oxHVyqpYAeMn6
MYLQz+x+bmlnN3XXuG6z3w5fT3Z+fP1HZCMhpK6ijHqUzYvAxC4b7+Sb6ICM0zZj7vq5gzu5uEMN
WXJ6lJOesZMT8wFv2jHvJ6TEFOieFqyMEpUx18/DIuxTzTU3fSCnEXPQDa0X2f3icVxGFw6icrwF
hApOZYPHNoLW/r12MLSdLeJtbp+/T2TLm06BUhxV6av1ub+Lkk60xLwOC+lRgNDk7qihWQTR400G
saGt0Xt3KU1YRhCZohJUzR7XmlDZW/MO92LNJIeYC+uY1CWGa3ZFbVR/28/pdno3Dz4H4tVRzOuu
2OR+wgGiVLY/z9KkLZ0OOm4HlMnGY3Hts79u1sTGXlbqjcB8JAcLLxFh4slkGCCSePgLiMRgm2lX
Ms3QEtIbvNz8PUY3vMernYHecS37AdqfoMWRulJKLiOidM2ofX6mJwxQJ8Q79AMA+ChoskkvgEeg
4B6XwrXfkx0SPu7/ik2ktv9n2+OYph5xSKSqyEVRFFF9N1YFfNy82TVkWNc8VTL9S6rjbyY3znvZ
9tuVJrsDD6oxcXAFlYsGdEt6kW/o9aRPN4EYYG/Evpa+132fjx4/ixx/Feo/cspV9pFy+FqKGNlg
wPUKdq/CZaESqzpVNSEO4MhBffbSgrlTndkEueXCrUJIEZW2g8DZugQvRnk7AnJrItwR3RIOrib/
jjZrCMu4jmCX8PH4wZOsP/tSIRe7wr4ej4o02aY377a5dNIaBLIPSV1J1CVangJi5JBvSpaqSLpi
e6QqaS67L42emCaKpkMhoHPlQiqoorfp1n5XGHZUwuE5oxw/p0sg2mKqsMvv7sJeolNC0i+9qkvG
4RkjCBfdnvwUmw2sxpTNH5uAQJPacfE5Hb9c+qAql9n/OcFO9+g32bCDp38rR46dmSiqGO2uCXTT
KsCsoyCCVojMXlK7vaRQeYyuYsAsP0Zdroog3IUFeNi30x+e+hvRJBYHYlYM60gAuOgZjfU+a05H
vdssPCjGN6IXL+eXzs9VjDAJmZ4AWOIC2E6/Zr7fy3A7hpY6Z5CqUdjCc3WnfWAGFmYNvlJON5Li
wyw4sE/jayDbLOdm7btrk8v5fmAO5w1U/o6Hy55JbkuajOZ6EjHNqnZlID8KLxHv9ty06E8hJEMc
UO1F5sZQpuRs7qDG/KvotczogJSorAimSfvrYIqCnTQgSS8nG/ZbgphTZyj6PxCTI4V8WI1/dPKC
yox7xMWcO51ieZ4p/cXp39HqOEifiB8SswuagfijQey992v2upSy85BrZnGIivwbIJS5V0J3hUAk
9q4KudrS61kYoY8dGk/dvcgwswmDx57+c3oAX+En6Kd5cxBLw1jyNAlhFJP6XrHRD3cW3vZLe9eX
blXQZlpDPBP7zaBs9Qb01PypxH3bycAyWcFHDOQUplNhhbLQTdeVjKX4NVQjKFnTV7GaclFRfbbM
aAsb+8YAhXPAFlYtQGz52p/IkOqWX3FtiDTO3s7FCH14ezgzEDLebw9cE1ZXes8rNAPSe0CKZS90
MvoYiSpE8bNLgQPW/Wn5ZHZ9RVaqpL6iSRccNA2i2PAlyjl8lboHLfKSPTeKWiymtA9enTjKLtA0
8Rmp+KHqEdGCeVGJAN2vfojIeFVzIpq9pJnAh8rJWJl/nc5DpHRWn++W6l4QTrBqBssg2EIWiDWf
9NhOZSnQz9JdGugnwoSLpr+ZMArVBlxDycZTLSAsfIYPPHVrPLXQpO7sdlsiutZhBFtvZo95/Ycj
qqEnBI92RXyixJ6FlwzO8lasTtmxJfRkY5A5SkawXI4wH1ICLGoa6CFKwfHlk3QYei3OPCWffKX+
BOAKX6MGuMdknJu2bwLjKBQwbQZ0BxqbObwOzB+NOl88BBGHQeMoyODmyqOv5qsX1StmsL9BLYSr
pbx6FBuzJlU4WkQTLbHbE/fFZ5VMs32Oavup8++lxU/dthbxlBJCTwuZmDYrnv640cSNXQ3uwR/F
BkO8Z4b4VW0XeHLnC+Qy/MLS6vaHy24RCym6f9hpiJvTivB6TrHZqzR+oOJu6MvwC2OnJwim9HWq
QD/yatitcjWdqU5i7om99+qORGIvJGOqTDNOetpDBwkBhIDs6BFKYNScBDJ7q8B/mtnp+hi3veUp
bppoYVfuDYpaJ5vwalxeY5HGF52cX2uECrQ0NuxjEcbCdn9RdgtXrXDKe1SK2mlnw3iy+fRUkzB2
aWOKKlSXtjrJzfab7ymlwYMLc+Gdt0pDmL/pEZRM4/5/sXewSC2gOMAv+REJivi5gNbj8BWgMf0c
KFFEtCtlLxx/Rs7KVYp4vQuaiLZqinyMX9bNoQpCZD6FjdSU4X6fSAQ5UKRRytTFriX8nth+bHPj
n32AkK34lBGy4B8UUiTarHmSc6Q4WYPtmy+e3U16mZa0UWKAyBbQDtptxCs/aN1ORQJjpCmuEmWo
tiI/+S/g/xscm3n5zF4idMcXHRFnEnp2bVJDLGibOjsJsPWTWX7M4OJ6dqKoJhrjAlBYxrQDNXfC
Dc9jcMqrDAG2WE1kokzt5ZAc8KUhqPO3HSBEP7VUhm452K6jAuP/h3zZn7Y1g/4+FnalLRi/9SqE
E7T8pqVvGZXldVI7QIHeNUGb3IE2Lhk9mspP/uIhTOLHAmjbdrYtQ/K1/7CZNeqMuEm3cdF0C1ol
NnJS2ZcUV33ue77hAZg2659pKo6cO3oCRbD7lgh1JLOdMgHPoatRJpDu8M9obPwH8EBtfrvMpQ4N
Rb+mOtf5ItJxlCe7pXDzPNfh01EveWS6pNQYxHAPVaqvI1omuI+E+2fc1EeJ2iLOfcRdIIrFBMLn
mruEMTDaLHKjMGyikGstKVKNCggx02Ku8kfI9TCxfut8ebW1WcJDDCpClgntBiTyR8+uXfssN0QL
KPI4gM5IaZIQaXeVKJXbs32uSKGuxVf5we2NwEfPigrrNepQ/E5UAC5X24pCPXTBw2WCelIx8rhu
uq/UnQ9K3R8rpCYPFxvdn2ELIRImc2hneBW7UyNrq6OfRS1TYgUTEaC3ByUFo3gr9c274xB1uoc6
YpJmpZiWIKR66BdpEYowaZuSS3XfrWpMMDRFhApgYO3f085nODDzCj87XLqwmLSB9vBQV9/fjtMR
bNLIWEaMLEG6jr+po5zP6uNRC1WAbV8a1m4IkjKnlXUpzHj5sMDHOXv1QQTkVWShvsbdpHtu/vfz
Zvo9FaKmI+UVw7Nkm/bKAhdltxSaBfIPwL1XZYnJJPLgv6ERhdReT3GsQypfxJkzE+CuZF5LKx+O
7no5WLEf0tMJzN1pEG9NHL4t8koyYeKcdZGjVFMsODjqXAZknOAM/fwTGejIwZJnyUVyED+EIK1t
Pcvm7oxzJFWBnVoptb0yBH7eZ+mOVgPvLSvTsRSTGLko0O1T7kO4dfooE7E7/sAmLOX/f5LBaU3S
S7CFkzQ45Z2rsKXoM8YF+TxXa5xfZCTdHJUBqCplrAL5zeL68TCgeWxh5AQeIl3iy6aNVi+6F1Ib
yRTQN+hAy3bCT/CMxiEPZ0MBBiWCtMl56B+3NWW9d0C55qFF5/2Dud92cq1VGGrPbQXdoWWhnIOe
R8qhUxg69znKLonFVygYxa3ySdgDRypiF74ckVb841pZgYSQB60TzZF8KMNGqSaXrdUMT+VAo6Ru
TmIxP9NqA2kHlanHe39LeN1O0wDc/iQomBkud+gwANLYCXLDzSUsIlcC3HJQIZXrX0cXNYDwe1wx
hEu7/rfwHcQdxZIoaCI2PD0P/PoSd2MVkVIkPrbs7+SjQ+UHn7ccjpkwCoycfyJv/5b5NR5CWwc7
dGYdLnA5ZyR4RDBOOi96arcaXRclphl8xZZleuEpe0JJ9NDLZOJneYzNeyZUwi2HPp2JUJZ104UA
5dlahzjRDoOwt32i7mUzVlP1mC4w57pGGsPkM8SrWMbIMSNCvCRFbaM/2bXlzUR8KYQuo5SRYvgr
U19aWGbu9Am7OSB7KrtGyC/S2O8GY4dU0+fIAwmJKwl+5DSK1rJcvgWcyluIUTWsXskCReDPvzWb
53vN/cPRz+PzTepIBY47HAzJbsjwD9UmcWRwiHbg65DrtpAb1DgU/rtRtj3smWpMRw/1BiaXW921
8diBFRxoT38bk0XSlBxTGH3LB/cvf/WxQUvluj91PSWE72M90wx2bpdlKTQvhs1y6Z2ONlQj3TfM
z4b2g6tJq22UXbEvcnDka/wJs8tbroWGjU/+iVaHwSP8kCVIe4nG3zj49wUYmSHkyrjF7flFj4Nd
5PeSSq1jsK7yWZJ1QrESg8z5QvsHrQetlOa/EmFox80KHc0yaaRT7ju9+CTNphlbEZ6hrCdZuDuK
i3QZqp3aMQjcyyHNYNcZ0Snlbug90AfBpOK+4M/NCFVVH/NeTEzt2f3TMtkprP+Fhspw9IIy9rR0
hZp3nTEE7wGSUuxdPkUl1kQGbqZOBAn8ZHv9ug+vQVARWVm59FIVTDe7O7qc7tlt8PjvIfFZjFJO
k112u4KC7rRhDrsyUXJWQ0bvSfIA7vlXyN+rtZSHdUnb3PVyzSp4HzQxuE3UAYaH74xpGDmzyoAt
tkbnG/GivToNv41myNaxAMFlFC5YuFTztPHnKYCYMZf0EnnXE+J9eLzBFu/qNz5qq3DGUOc3Cwxv
qXtZTvwu65pDzrMJVYnmZ+gP8BLE/m0NNuEHb+pkVREIzbPQgR/ALZLxlKvkaumCUsGjS0R8ULG/
6WsSTXu+8EsHKg+hy7ROYnd5Fg7rbFKmULWDHW7cVN7F/4jFwYn+Ea5RpzyRN93hfPyJvpAvuPUV
Ja68Mv4De5Q/VbrmQJtQ8XEYZc9XUW728WEE3f0834oVEbkRrWJNYgkYB1VG2nkMgdjxLC0P88Sd
9yfSr//G5+rJxpJ3OZ7rWCgHuIJNw2Cyl0gxeKM4eNtXCmbdinrcVcBVRTnz2kcIVHy8O7HqewbB
PDnB0sxkang+fo/diaLJ/llfce5aeYrXnVDdQ6FtW09k/oBQqpuZsKs+RxC5D1fVpEqiVr8iBXuU
FK8Rb0gHKoMi18XaP6pwwd/Dx+9tX7MKNEZ5Hl+ZxDnSbxqAODX28KxEZKNR7vBYyGFFeiY7AWjF
FxZAC1z5IxFaITwG/x9p7NiG1TCQ+Gz7FDEN6GidP6LXjKCgP4gKnSOq3Ws3prN88o4LlKbMRWkw
9elABmSGbW5xaOA8AFQRHaVwnv5DTQuD5zMljO60upDX+qBBOD6ab1eIDO9cKe7c2iVlCF3IbsW0
J69VUvyw7pq6RgSiQ6Zf9cOGpKDQJvqSSIVnSVBIsXE5DI7a6ggRyV9XN83tZoHC6P6rkNySlvM0
F1D/s2FcEIzvHFwYTdoEesISRO2cj4I/FP8nQF3apGkTL3ehrPWI+aZihFGeUyjIcS1qX+zbYnNz
i27pA/J4LoP636anNGggQy0wLDl27a/Rzp/r4wEzq8cc7y+RVdO0mzZQ5Biw81HytBmrleuOnk/v
Tt65WanSOcbmj4bFZAc6JnqZ30R2pkxMgrWyBVS7tc/+FdTD1Dla/HJAdd6tmXyX0A3N87TXboIb
HBkFpJGvPJEITqLbO9ANuOQZbzBP7DpkS4fl1Ct3uCk2529/AAl8bp/cI4e0NLSzssYltDItbhe8
xUOratPOh719fnm+sgL27F37cjfAPm18hS/4fqgGoHKYrjpKFlaSm8MsytrwtWp7ATn/hKEVZe4t
VmuQLsImqHx8uNT9eTPEoNdFuv7HssVLYT+rADRsFh2F2PozmRw4fotqtk0Mlq5yMEvdnPqVWQ55
PCvg9ujacNP13Z5MKYDQMDAMZhWLAOk1c6IuRVG7tgS/WvJy5j3sjlXDny6eBFDdf1YLiyitcOSi
1j1AnOPU889g3mJi0IrVVS4XEi8nT6TxOlENsdPpgCrY+APZyAUQlYsY7VzujZir9yPWvhoTS7Am
46sCzPdL7c5nb4OkYSKxgKEWgXUoTUkEFepJMqZuWZxJf/tyeDgnN/mpNrUJxQ+KQ1t5+58gUtKW
5POKUWiFuP7u/HV3waWjZr7RjQ6ARAz7sWC/71incqTDuk8R/0Yo/A36aCESfv7BuMWFlGk6DUW5
iFX+NOfnlK1cEWms5LwZFH7Z80c8q6rB9oUwrESu6j7UYYU7QkOAWl308wAoQwJY3SlhQWnn5lS9
FloIdGEtfqC+FWReua28CDsdcraZIrRJi5z6YU13XY6wtafsy0GTpXlY7X9z6o7sPx+qqgSymPwe
Mp4jwUlpO4E3GmK0PTRS0lv2ewktAt/cGofX9ZQ4bOl+ujbCwiYOE2IynkDsKmOtw8L5EqGe4u57
KC+pNkn5rYquvwAmB8oB3qFbo2p+64dEWs8lJ4/IgydZnraHWLbck0pUyPawhJjeEs+JWEbBJb5O
fV4KiJ6y57Cwn4/BVCRXlIsppQcGVyDJk1dRd0rp/w9AEFN+zuRZH+KnN4Mfqea0yAOhcgxH7o31
VaWQhK5pisc79LNQAclxJ38t1SgWByJEKsOJfqLIoY5LUg5xXV/vc5fAb4IlZ2RoKYqIRksv32OK
iQ1qnrgqi+xbwjRFElhs2c10OqcnNakBZMWq06hqsL3qRTnYoOwjxtl3amh6qtwaMcFx1D98bmb4
fk8X+GX0W1PRpjIeQwfs52XXkULOemKOxfzKbi88HCnrpS28KMnuD17lpnorlUsoiORnyu7Taswz
15FvglHXgNm4VPrLpydLR+0RRavSSm8w92c9qGmADQn7L3DOyDWQwslFEuanq4f1wyy9J1dCuJUV
usVXlZ2SOALtQT2x8zs/kf54u10PWKqMfrGX82x0WXldg/Csqk0QhFCiGb61EKftcgxDCPUzUNeq
/z7DsEDlYIah4dngqsX+3ysLtq/3V1AZV4mjLZhyedIhlVSVI5GPuQLwYlrKt+AU8DLJSH9wdMrA
k6Yry/KXIKQ7G2KqZ++7BbLnON91s08qNe8vkhrfKokmSZbM4rip1XJTIs2Eronl8q7xsfQ5+e1u
4XmYA3WigHupLtl7l2klyoaj8C3f75U9cE2de4sR9Ahq53KITjI/Mb3zZ2jgnv+ixtrJlmFgn65/
aElF2Q6gmzIzuWcdxfRXygmg7ZLhoyQhZH9aosz8r7rB95VH4z4bC5U/ZwLE+UBRO3UOKGaNqm8I
QTIkBB+6myhMKfDw4KNuIpNWjUXAI3WwvJw7dqvMDUJrKhEf90tqvLA0Judf11NVHHoJWEP7rG41
DInMwfOONIn4ZB8mGMfXCByXRD8tz7UF0Zht8MYZV1KbCA6hXMu5jULicl61gNoo59GrC8nmN6Qc
8hNDprv/m+GnBwnb6YtR+uXW9eb8Rm11SlqQb7BkX5VyKMKVlkyZKS73+vkWbP255mKdZFwz1/G+
t3BUzzu/bbdN0bOB4A5sQBJEJ9SSm0EMRj4LPBGyMoElvaO5WeK0Zd/VLUbeMWTZWC4jMV9rkDiA
L732nEHbP4pnNMxNAiBWc8zmWnvLWcbJElQbeP0wNoKdQqTPUCyskaUHXzOmyECd+Ijk8q6R/c/K
uqwJg3JSBpJ6zLHPbMdhHLdQQ0uQj4vjIrv+GEVESs/PrLhjKnwDHpvuv9xjHFoW6oHCNp/mD47A
CI3I2sv4MNvzhe5AdI6bA8TqMJz4NSLF5xpv1kJkiX6+tdDioSnrpF8zHNBZigQuTvi7PRdcO4Or
btAL4RRNTZ7wLi7clxmMHf7CLcFTQAkfWkUS55mvbBwTrZfG94giWWc1r2CApXiqCO45XJ4X9bSC
zqId+UCWJ2EMzvVOteALJ4rWuELnR4MOQT4eujfVoXPONSyswaAaSsdExBFMkZXg2C2DJRXCqPz6
+t6EVNXjQYZ0+HhYX94tms5TQZp80MenYqctqd6ODGlddbF8DlIGvh4kYQ8DU3Vvw/QKXZ8SNAFe
vsi9Zu/bt61jjNTyWvXRZ41KY20tlFRFSm+9VksKVCpAFRM7oUsLM3U1W97kds1O6ERXfE7kJnir
Albc8w46D1iKzPHjxpZGWYYjYuz3UldCKFEzqTjoC7aC5bCNcQAKqvHEoBiQEhJBQD9dp48AZ2eN
Swag/R7FhVuA2XvrBsRjpo+FJb81pTBnPgINtc/gopmPbjqF+tEvGquSI8An7F6YL1AnahS1X6pw
v6iU6H48WTn8GPIInKgEtFRHHeMc8VWVIR2XZfrut+ZdAnCJAOSrl7mJDTjhla6ogyWTDdi30/ja
QoK/c8cJf8XK/Y5SCSe1aq5zALbJvgYAP9gmWPK8rAAMpIus5vjy74GCKcvjG6UbCD40NcSlzsvY
XPiA/aR6q9z9nBz0lGaTJ/bhJzb2CvWxL7ehG2dmUfOiEOz1QgBoiaqHIO5WgO5UbYVEqLsTtBFJ
VKFJ/jjhDM5l9rtzxB146CT3LGetfoo2FnthNeSkZDbgc3ldvzuduu//frVXP8Wrv7OX3GL+AqI1
elkhJ3A5fyxlJSnVAX8oPIf5eLRERn1hEtYiliySlfWkQWCTeMh+aH64sDeYc3OMhtjccqEqkOr8
1SEZEwHmNZKEEmCzLrC1NpdGngbTLMbM9Fflp13nmdMrx1is5/Sb2uMgKCHgDJNLyQEoQGWsL5NA
/Z8ZMqwn+oCqM8msdbE/xoQVa7vsx8eVtrA8TB6el99mrx2DsWVtOKSQ65aafAL4eNp/GS8Fze39
oTz0NTPXTcrwPXBH55QZZZ+S3GLD9NuRMLmbZzuHHHVP3SfBorfMZ3YzZ5OKB+U3nQLO0Zp7Sfh1
MCOSlg9at1IFiGOfzpBd+orceaKRSKrXlOvsmy+9hlvEYXGSBxr6uwu/dZy7GENwuh/sbflhqMJa
7N3jnjbeE8OdQfm5bUmQ9naaRJiC+ch7TH2SPPNshNmDU/BGRfDUQTzZWuJi1nw1/Do6TzJy58v/
2eSrTGi6ENbdAMpWXfHTgRRItDDzCP0p/Z75rkK8HyH9Uy489YW2eCKrp3JENPK2y1TUCKFKfy/7
F8cRDJBEJwv+67syYVusQ6TkfJRBsChPLhEn5smlRI8/KL5wXdQ+sJ4FTDW1IKRfurHWrUFgDljJ
+K1Jd5oCwZovjihiG3gWZJpSr1CZ2C0nm0kbxts/hFyG4xSgMSR8avL8SzlHPdUC2VI6AvmV+vFN
dtwuopdfZF5qgxdMlQRgYQGQQcQbimKWxEHRBajlsTnecRrsKRR4MNNBAOSZ9M4axGI7n+tVB4EY
2GyBrW/mv1t3DppnNx7a6tUL9RtRjcYqfLJh9WBAUSSuRtDRcUkiERJX/A9wsUlz8jk6bqwRGYyc
ZNPHs/jfVHeuKn8tkfEVlQFmOgt5bLKLuIt9vt5/dRPLDHHAhPUdIWuHNrXz9iAwvF0UEIa+ipTC
iYZ5ysiSAXS2vNl1DuLMZQw2TqjnfpUJqNkOTS2pgOf0SUm8vaSxhh87aRPJiOkUnn854FdIMwMy
DZ5AQ8R4s1TRPqGHm+blMel3gbI8ujuPHX7Z55TlXe0Z8ZwK1phWcAzoawpAaY3Is9CpWxaEQ+2y
13Wiu3KaTtxt9wlTTsGIcZw5sD3v66z2/dPrq9tKuowWUYcOXyN+mlBocffCK0zrjLTiKzx1u7uz
T2kWneN2OMYy1CzlypA1J0uNjpo46BzyI9yb7KakhK4GamzZy0zMDFvucbBXVt+SGtWj6TYy/8Xj
1IZpn3wuSqn0/U2nxZW8ryYX6lveHjOVYBOkcK3Jx88vvm+8sy8nTq8tUY1Zjqb7Ct+q+jfrwVED
NsijvPTjVoJxi+flxUbXKQcU5amTPcBH2uiDmgov1OFT6rjHrOf6gT5u1xxMYHv40eon/GuiqB3+
y3CrjW07Cr7kLI8wJscsILueVRTXMUHfDCAUTXaLBFTq0f0Zrvocr2NNpYv0VzSAkRAHkg1AlOnD
7GXRfVyRPsNj7zAfjfcaNsEeWcFu2o3lNC70uEydyjG52IpiTjMYs4xRudjG5m9wSLbZdgYBiYcb
pAxCcZ+D72x36gOc5uoE3n4iFJDmWT6pkw6o9+aJVXpYinLwSndEBhcJvWpO+YdOTyhYvuwkprSs
nb2NgALZSu3r/Xx1T2XZ2KA3iMzSqMkKe+DRTnkP9CJXEQPqrXW59kP9E1aiuW/xs89M/OqjtZfu
uXUB4qyut3LqfRo+pCKWtYET/f9d42v/XOU3s80r4DLvsBKzF7/SPb2PDY//FpfZuuZ92Vfcqo/i
jQ4hQUk+cy/8qHBUAAFEfovwiDjQGLXVCiLxX1CuYYRCDYxZMjuBpgMqXKtEvykcObLtWnhYVMH2
3eAwWOWo+31A3p8+x3g/PyY58VEtXMwa/LlSwFHrBjEA3PoB1DoCeyuKzwrzNn9olBH/izXhi581
PBeTXDK9gOPIJHS5ZZM0R8yMGOYuICxqwAvbHkso+HXVoHLwnIN88Zb05ClUYH23AKn1cEeb+tj0
DR+ExMZCDdKtDSWWHkGGHLpc91dFosWeeOEsbNlFYTwWngX7vdMb6LrgoyOkjoUDOtiWW2CVHx11
hEYHpWA/Pl1MAPSWhtNgmE5lOGWk0S3nFEY9uXsg2QqXPz9o2zoLXRj7CWggJ0iY0uduTWFQzhTz
DNUbDFNd7FpL1RZB/HiDrXfQ1LAtE5wO0Z3UMABPSesdMze2cCBYgleIi7wz2zY11o/V68N4yk7u
TP1Li1XG3btv5VBTzxxcPI9ukHIyE4Ap32YhHwP3RWFwD/A18KW+edRejHJQPpEIP2MLhVSWcMBz
r2gxYNCgc8mUc8sasSamELhCCqC8Tk7Ae/1YbVQLw5Jwt48jRLzSksKmWDurPahjme4bqWN9NRNd
zQo5YVUgmeISPUeAnRR7Xi6jz+o8Q6+aU7zlSVyHw508o4aVr4dKHURcLGSM4mVKkwGIFr7dmdwH
ROgrpRxwTytUaOD0oYOEfxlCp0a3RaEgK2hI2kGLgF+vVSKbII43fj0tVEo8daTSKneV8x+e8IQj
zPYUR3E4Mx7PbwBER84ES3hLZKwnfxtwx4mt0zXPad48TidjaJXdOTm6i5EN17dh8+RYolt0ijSe
1O92rHRD5fJlqun+2wg/EMkZsY42/CihS+vMACbF4GMFjTnyzQmN7SQwoEgWYsEXa9TW9uH8iDVC
5ufjmJqmL5sc2fzvsGH5w7gFI9m/7i+k1R8IlPm0i4Kjm1goaw92vmqhT07ca/S49sEsYCC1zW2/
aDGA9gwFaElWhMJxbAixbLxZ49nxUczy5jyURd27A3KkkLoEum85LFZDvTl4t9yYSREyvgqdTaFu
2vQ6cGd8L8P9Nu8anDrQt7rxZa1KuUu4LHWMmCrfKnGkb0rCueC1kIMpRk4Xtdr6pEn0opyqOk5G
BdtLxmKFJ62q8OCxkyWE+laxibWOXvj4+yQEoA2s8fkcYNQTWSauYQTwqWhuIlZdSlAdWucSsBZe
DDjzFWpmuYVOwRaEKA+jtZSc6aatlcSBs66/RsNbmTSvi+YD50wTqXu5D2gVh5Yi+KBoU3IrehDc
OEpS+EW5vbzMTpU4JE4qPEKfBJrxtJJ8EDRGZJHH0o6f/WfNjEhAV4YYkIatL+qRHJ+0prQT7HkX
X3+2/ByjW0X+k7dMACS2xpV07OamyKcJsOij7n4qd0OzINU8V3+iaXJhRV8YdWGIAVZKtqVhw6Qo
ztjFeMMKLSrLhSh0gx+NBXQhzHTHU3XxplTjpMjyszNqPiuSD6XgVmy+qSJKmbPUczww/qzI2i4X
QhWMWL4y6WAcffjUT57kjMtgnkVeQHmriblY8lkrsmfBgdzLsSCjcmvYd2dh3dlRLlRRozZoniAI
m1nZgMyVTeMAbPtnFZIdQ5FOcVP8ZjbRU2OjbxQGbTybS4fp2T6/ND+9R9Q5cSSd+0WWZwxsJpBk
X4Z4GT7ai7WDkuTwWa79QfYpTjt6f9G+ketBl8cOHxl8uUFtfnczVamUWYL/3XZ/+r2DOlJ+0b1o
TMpVckcsLMtv3lCUZSUHHCxG/abm2tE8veYYj9LAPBvlKaYBShQ8joYrXhpe2M4x0hHH7ecPJrIK
qh8kZnBodABqCvmocGpGzZUokRQKiOQ9k7k5CEqtcIZNF8NiVuovj2W+tYpl4ilXqROCkBW1oHgK
3ywCh2GSrqoIJ7yOqDlqOpqytIQtmw9Wm5et6Wd0a62ShPTDTnczFv96J731fXwgmwQZDI9jsma7
JqNw1zr273k7r00xYZ2aN7KyC4vhCJpytwBMOJUc5rWFDpcOmAOCYoQwW77vz4dl4yw8AKYUgmAr
Ey2eKcTlRNYODsOStxaX3nnv+EA7x8qu7QfYu2vT9K0czYzKvxjXgFjRULMOnxSTqZqGfe9Tb0uq
Pu6keEgiCmK7DRmA8Hpn+/8Byshum6tOGNoPSr7XFlh7q725DbCXlEUlKizYjhsA6CFja+5OUROM
S/F1a9xKrod6VE5l7lGLDB38o8lHHqorsCbrj14qT9u0XmWOFUwinGeiVYXwk1cDOBsc69xQqaOU
4MvETdJeJPvvMp436ZX87/Y+Aklg34N8qVhOR2+kYN2hux2TPpXHZHkjjBvXToiiDWL9IfMIujQ/
Fn55/F+gYvYEBhbSlSMMf9WOf7AE4FAiOxZGku1VtldvLK+w6tdF1Zm0H4NHg+zVdqZnop6gVJTJ
5oHMe/UJVDlbtcyt9xdkFK5sW88EvePkI2MUi9G6+qIZ0GO4NA81ZhI+IidPmU6g3NTp+5OED5fD
3kSSy9GOJlZ/faovZ3sA1gci9+Qen7Z355vyz6BPN9eCDHIO3nzZP/cZX9j4vniB3lTYSbX2ri7T
QEwWNA48CiChjlTrfypEKU4ImxrWgLje1bUKOtv03n0YEcs0rcopW5dJ8Xhq3ONUW9lGPEymUmTg
6I+3sBlLHmkw9Gfyh6w0re+YuPjYTM7vIW4TqQpAfIf0nK6N52iFdkj9kf12zgqSnLH4esyyfUK/
4DSIaD3PAqxAFFT0WtK16I/BBzG6BMSXwoNMSaeBnQvkFlX4x1bmawn5J2k0Mjr98kFijb6ghbs+
/cXWw9UsfzxniJupw7jobVRL8ITEOFM8ruyaPBM/crdmeT2zbj0sotSSPJW1kfwkqKnyg7W/whC4
heyM30jfYciqKW82vthkKp8b6k6E+iMxMTEfRqQsJM/d4zn4+Ueke4DmcdoUPEHy7kqjjbT68pOZ
dg9XUMMvWvgIh6H4OfZ+R5q08kB/xoiAyGcAsNiszqVB9x863k24gl/FCrZsssbiGpPbVaPgu2GY
4SlP8v3jZELNJMdrc3yHETj0NTAmsFrLt6RMv0iBqF/e57WRSa6lyVT3swdpIduwyS1QPN4xNAVv
brky3ZPE1skUUF98ijjCXrKKapPpyJs7aqldH4Ez2jIpiz3FRk8wSubDw0CbKYLNlPU2/U7QF5e7
Whd7uigITFS3i+XuPCNUO1XNXJ+zx90JX4VcwA9lyLL+lmRK67879b/CZbujRumLcUtmQ/97Dzfv
K9+4tfg1SCmhJaVdksHOvKEs4vkSMAQklcQlJDGiUJUF+RXIt10TFsrz4n7j/ILN6DorvNetLQWb
lbJVoQoT7j+Op3IFTt3d+X65lsy6hfhbNsDijalD7yP7XwbzvABeLVllKc+Gy6X7AFhVzNK2Aryf
pKZpYDNkHa/U8Lwb3m9m25WlRzPSNB61ubVYI+Qe2IuExj89GYNGwIIIQ5nesj0MXYLA34Nol6us
o/+xIfzytbhKnXhChqM/JY/VJzZ0p4wFDn6ge0Wfb9NnQS2RhS7UP8X/E7i43wMDAghiczCRMq/K
RdJ/7pvlfcbjxVumtG53uq1OqHkRw3p0A0SCgThs+4FBSCmqfAHl3zxYyLgW9n3TCuxQs/AIEN83
gJ1fsL7s8RR/Taa975mLrmWGNk1S2BNYxlHBwSpMLNiC4TK/SCt7IfxkYYqJJM4IYjy34JxSkg4P
S25xKbTPKfdVw7dVJkS2z34EgIFnwod71jl384bumwLAk53rVwyhQb2eiLR5MiLEvL4PHKdwOSQG
w28v1RQa3BkIC4OrVJpIRbTsTK4Opu6nHH0Xbnrm1xvw5hLZ550PL8JrWPt4/ATxiEhdlQSp2XtM
PDdxvt858vSYBkCf/z1kLO3wlsEWvm0ObAdwWXvXTehFlasEVN9b2FSLDEn0R3IsUeJG5jv4APt/
afYgWSoLFWmdY2UbC7om0o8sOH70Lshjk9G52PmmqJrUMMc8kNB/+faVtCiyARKxI/3trTkKjL5Z
Vw2MabKW58gR6fQL7plFl03aAX3uRxHo4eMpeRYYOhikJpbxAWzOaHPwFvA8A+kEV3mt06DfUV8C
qAogGP8GHdABXgUqzJ3Zokj9Nkc4koebCIUj5EgzpNFXaR7/fnnXKHRoCOCBdSPNsEoGY4uPJzk0
BvCqj7cQsbAhTz9M7jsf8JDrdtTajbyc5fofGlSfbz0rsxvDtr+DDj2GJNK9F7JL4e1AuPvyHdem
PXNhDlVitfvKsj/FutIQPr7z0un79H65Cw+Xng/Ks3JfPaTsd3IK6y3zO1jaFOjsh7dr1tg5u2un
UDjFGVwbjRxWQwHevZQSxekUhxSt3nWTsBOKWkFU2FHsEdyPjUW+HQn+LPt+5OKM1d/6LZ2/zT53
NGuxtN+XLdVO0Ti+zQKpghcPOg+yKG16r1v9KWeuk0/KtDNO9Zfu21yH+6ezoof8opQ3MO5hPsR1
wcDIviRmLthoIFxcYmYDBniuzeyT+lldcNY4UAlRF8DyZDYLxmsdlDD8sBXQdCQFC2JjBQaWQKrc
Z0pd7dyk/nPPf3iK59iWrW/R66uVgxt/WY+9rrAR+Qf8+w0gj/Az7iBKmgrNCn5n02GLYwzSM4Dl
oRmEDictvthUf1OcNSV/dc5oH4cJd5VFwb7Ro1VO0ji3jemn54yOo3iPG4mbTficP54sdJ7ouFep
dScxXl6fixwC8nhGQzJ9SFPfSPiaUSLP6xnRLKdBwXtG1TfSz+x7ZpkmXwKb01OonzVhEUvj8GFv
Nnpllhc/To32ZgU+QFuWigZLTgzxMJcp7iMzky9PxGMmelRq5n0dZSDViefsMqxEe4g1yYC0aHi5
WsmSRcisy+SU7E/1yRtiKMzyuLxk2X/pDo0ulrQ8gzuIm9fjGPvaWe9jfDWeF6jikmvlDcl+zBZJ
w9aM3kpQ0e3C12DHWi1H+wxVkYR1p6br7G5R7I/mFe5O01kQFTirTGHB5Uq4cZEdgR644pZQHA9W
zV98Ya9FPcIdY3weNdwbP4k2W0HP4IY709gQ/9aS2MHVwaaAGoiXupbKUqifoOYwlsF6CaklNTcl
LPgU7bRouiYdFgIQEsedhV7GuaDTL9+Lcfnshqu2iRz8KgMYHqwJMc7T1qMdi4xjGkIKTiZi7Uw4
iXbRt3tMoXY2GN8OeX7+5bll6wcwnugoej4ntmNOeLCiT3waEvFNz/q151XOTdEb7+CxHn5lXF6E
DDpFqXYf4MFMysPQsPbXBCK8rxEFAmX8cUab6xQwYOfKZgXJV64gjtr6tE8sPOdqq9ha2brTFtZt
7kiQg9+lWwhXXItmF5LqVnBQS3nKY3nvQqXuA32bBtnuArms+G5El4HQQtnrD9TDgPV77eS7wFV4
B0gnZGMTbe7gOcQ/J+QtmO8FU54P3Bf79eKFEEmHXoc4Ko7cLduC2k84HKL0gwzmH6VM5CmvvCq8
uvgmTj+XFcxz0ZO/a047ZX+su7aq6aMMf5y/pU7EG9zySLTTsM5QnU/fmz8H+TjWbhzMGTqcTgLv
KCSufg62DcFciMz1A1GkrSyJVZ8Y6oh9us689147B4KNeRVvg65Q2rfkeiWPSTW67vN/vMmWOe4O
Bsyn1/yJTC7MwnecdsA8H8eXOftxz6up+FF5hilqTNoHZln6e9FrNhZTiJ9ox4S0kADWBJB2Bfi9
HCqlKjRZz9NNRUitAuxGGCwOtU50rbC8dAIvAkKOs3LLdZ98PjTEYFvwUC/HLOVH7s1D5Nhtw+ci
cvOMYB3ACfKei5RaMX9dawwp+uYQKUvE+j1g4Q34jc+LRVQVeeewB+JMwsbTbFvQKE7Q1HJtI0DQ
7kWXGhtxKZ+cYxwlW03jhOXCljFsWmspMQKSVKe/qRLhHuvjfavrvf3IAFeWMdbQ6H9DwP/quFo3
EKQAQNJbOygVwQE5OdK4K3iH7N0wsw+9obCKIbSWaZL5W2ClUYBcF8R3nHGT6dNsO3doSPYsk7iK
SNT5zgYS04ZqVOhk9m0BDPFxk9rDoRn1bXxBrkOiILrW/k8Kgyaomvet+x0Bg9tnP3WxzV7GoNOJ
JN+xqg4+ULtRweFrKX6ZGaU8w40B7Lhj9VdITUrsdIH3P3rmUXTf3wRUuXU6j3d8vyDzTynPRDfP
Xaaz6PjFtfhouYsjwdHFKWoCyKekUiqebD+steha36MrjRzwBe+A9J11ZF0A1pcSWVzvqR66cW24
oW5nCcX6hfJORzw+LEhadu+6ysPwtIAP1QD+MUzHs5C7yvMOef377ChJTCYOzLGYTpOzDa539M9+
PNZ5i/zkoyXSXgGHn2pp5voDjtYVRuxg5h2ArlQn+5nYCd0TfsBMmx+YfykbGSNWZMrcwSFg7RZu
fF1Gr2IyoaYMYSLZOmV/QsKO/gBRhWGzN6LAh4uYBJFuevtx+ymMSXoKVy5C3X5af/gTDhfnuJ/f
KnWDyewjVORQc9gTig/wnFuJV4RxHuEvs1F9RyAI6FT6TEGoVGbAP4KO3nvQN8cmJVXq/hi0cS47
1C8tWwUS99nv70AkMH9AI0pss0to/eAljn4YP1jB9PXT3ie+DwH/cDVzF85MvpM/8+XoqMng3Byt
3t8abG6agmmG2EK11lPtKgiM3DWBYWODNFiLHMDTvzHitYKfARIWA+/PozZhHLBxDoyAGSkCDf3t
hfP4DoIlFQWAOi1R3AbpCDeU5E41xjtmTLJy2fUASCh5QTyAJqXCzIJbnj3vcENu66mSQvEtlh0c
TmU/K4jTmwK573K6zVJB6KZ+LqYQPuzGwEJW4bgMySdg4QXGj4ZEMtjGayaWF4ME3TEJrGwl/zdY
WdcFDd16mBfaSZEtXQU0POn89DXMqDyELMbn9q0ElEVj21SXZ2msHrQEG4wqiNUCaACIgwLlI9JY
jlljFV/f56EtkMj5tNFoCzEhhhCH4UDXAcCXWhHdg5cU9NN4Ab8U+qjAZf09VrWp/3ksKfZpOqMA
puoWWSZ/hrSVZgp5a6Gi4ossRIkqFqgJc/LYXcBo4Ja2JI6A0cUvlRUbMJtfV+dELKRtNuqxTqW0
7SlN+fJL0PQBsZrkp/8KQy/lpIn9Urqc82abXAKv4KspyQQ4FbgKrD2NgPx8vtBwhS7L99nRbPsb
C0RcZ0EzaulyerOAhHmbWOEFRIVLSFrQliXUJh/0haToYJ8Mf2pRNgNwTYcbmg1T9+hilbP+VrMg
D+MlVUt7CW1UqhjqfFLH5BLv9BHEl+H90ruhTw6WB5dsOK+QUyJcJPdfh0YwFhf3QFCOvl93jwkW
C4Bi/Lvsju/2Jmo6XEuNbjvXmAwv9ac+V9uIWzCb5UBNOApm/5gUTiQUVzuf9L2Ev712nxLRhZcF
egDzjwrZ7/Y4z3XbNNriMfmdCwumDsQLrtCjmm/LlKPRn9J2ujciJJ8jHEjf1iR+zy9+TPPu9Oar
4KMuS9hlnrxp0ZjcZo5tDy1F6abSe2hL/PjJqTfPt/fWgDbH3lMY3AHzxVHGQO7VURRrZg+KrWav
r/X8HZ7/hLKxPXHJF3Z9WIysiGpytBS+tytqj6t5tcaygcOChq/8e2Ls/qjOr9Tq+hHTMqd2VsA4
crmfKliBlK4VtSld5S2i56OO14L8yamDOeZncKDGWPfjDLEAiB0XFVJ/cUg3rkHg5bMAlolJgJ1L
QuLgBgHsjygzgHKh+Sx9wJFbSm6zZUDSjxOmNIdhn4lfk/R/IiJqvVGKJMnqgvXDphm/izh5VFpn
SiLIFW0GYs36kMBjAugxPf/jVojqU4Q6QOch0MSEo1x8XH/R9JcS9LGiMiSX6gcy/uOiGVWsMfEA
Wx8gBzWdThBtehD/Dqwp6QSr4F+x8on9XBrSziciWg/sR7H4EVNctK5KPYPqNeYhut/sU7Fbl28P
X6H5uwfxE7h0AERzcEDd7kuegpzfgpfKEzNhocfYsuj+5Sp4eguBlRADI/P9FXzYy6YEOLs7cu3B
rSQUDnNqFRe0I3RK62Aswd3bO1HgH47WqOYr9MRkx4cZslab8gEEO+HhpmQ86OmOko3VMOOzdmQZ
7PNxU6NuZi3e3ru45/hr8szcEnxxkdZabzzXMhbJwUA6CG59aD6+lBrLzQ++J54w8BXCEYhblIqZ
BNmS1j4wUYS1YVK1BtJ5V1KsFuvJN2J+kz7gDpw0smxvClDQ9tuIGTKHm4K6ssaCl5U8efzOj9dh
xnR8+bXVPE/aFZUesb5Lf/eLQ7l70ld5wpcDPAxgmdmooLYy1X+ciBj7QEO65KrUX+cH+Js9DxIh
s9VvcdN0fEk6sGhUObQt2W0opFotxoxjisN+uwVSTmXDROco8BG+h9/YnBFAlbr2dgE8uFWvZwf3
r2oafvXQ6YySmsIyI2VvPWdCXJsUkUv+m/qlOoQiFYVpYG0k0qPD4Pt6kXBEW8Y+iYPBsFQ7ZIfK
68oa4Lmes1/RGLguNtHoMiUFRo92A6Nk1Ykmam+g/kmwFEHT71Ob461GKGGu9UZldwI8A9rJZ6by
Va9mEGipLJbrRdfQftF6/KyIwXf1SMv2MnkAYfKqdqwRQDIzqsH3syyA37PdwHSB06VSmiTffqew
/f7j67o/HtEFt6mw760QcHSvMBzQdPocRn5FmQYvVrrwCc+kncBXmLpDQQ/3rnlR9u69KGlqJsrd
x1EvYkDFvuAcSsif71m0PijDSnOJ2DerpuGyzijCE24t38Td2EGU74iOFUC6o67wOnbNfptqm08u
B5Hmi1gDxXKiqH5pzOtsxE3nymVPMULr2rppWzSv9ugZW8il1GaWvgU/bu34rIznVSR5KL79KqOV
RmCoasayBvypB0WCSBQnraaKb+IXyYz5i5ePzEmwczco06bRx8y2mQTdvNmIZt4lGq50E+NRAjSr
oXXnWt13ikYrd9LqkjR6ciRiqqsug5y85A73D0h10qYu9v2Khl1WzgI34mWyDg+QbTLTdsWnglq2
415WIfJbbQkWKQB7odz4zbhBWiErU8NHj1HoK+NO02rVwfRQBO3ovEMje36j/Atn+ZKpIxcHcyYW
vLRrSH+WbSOQjRn1fSvJCHAHARlQA4tvu977l28T+k2Xp8BpOEEbK6blcqFC2lKiGNq4ndui9JOj
dPmIcXQvgM3gM2gbPm/9JPC95Wy//8E3DWRUz+FG4RGOkwo8J3FvzsQ+BfR3oY0Tgv5+BTlNV3xu
z32aI438/fjAtuSyurIG1bStQrVmoREZ1XW3HA9VIky6kgRp6SEiJi+DanCtffHxx/EzHWZtSILx
u2YZb21f0rHyiwYkKMDVSmB1NqJShNh42Uvpze1FRZGfWAAkG19ooaTHgMCUhJRIcrMAs+nnylFf
6cA4PN7mt95HIgYq/lAaZKbHVn454RyaA0c84AZVLjVPThjXPNZ2UuQE9wuV1MxcKG9fIeTKYZOq
ZOCeMMrVT4U+soAHp+U1q+WpielWKb2An2mVlWMUuE3I+kn5cltHVslQeP54nNxZnJpGHLfpG4lo
8GiAeYkoCDpoDanfqEYUus/YaWeYjKjhOpx+pTA5GT7uko65v2A+tWQHIksDF9pXEKDvUNAt2AMQ
Gka4cW4SC19fnLPkPx4/BdD4TzJx3GIrktJoNM9U7ToxIJb8Tk5x8BoJjObyttb7oNm4QXhNuDTw
dBcMpMP8po/8Q2/ZKtctvDHARE2VqVQB+eAGxD8sPFLXkDsYjmYYxaqIBiANjwVgjF7qNb0yWr4v
lLUMJjNJDH/9UAEiYKHWRuvsQJJyaXODJs8lCGC5bL6BmPRwgPRyP68ZAaRLR/e5EgKjbSJvy1oK
epZJPjtdVXKCFodg3gZewzZsJwD6xHEGWA+qbvFVAhEohKvnWi5Y1KRYmE8kOzA1iGnILdlpvyLY
Bf/HfbmFWeJWBwwSUrLSejy1MgaXePtC0kXWT51k7OqumJKbGCZ8HCa/Q2EN4Z7vEmOG7GiOX3gH
bMWWSk8KWaMTHsq1yJkdVDThWUWigW6ytBt1riId3Y0Kp1qVL9m4L4opvRHlK0ZLmPYmKsSc73g6
0+PiJ5rvUCPhbgiH6VJldYH99bqtR/is60DQ5mO1IHnja1Q8f3wx7wPV/D7Wn0/lvpr3e1/HkquB
1wNNwgxDPh1qY6Cgb1BhwM+klFdsp1kzlTfvwrnhUN6mTKuQofA8Jx1IAAMDdbcfa2KU2F5yGfUH
q/xn/aMmzkh2GQjPk+ckqH60+EYtMjfD0kceNctlwZAptngPr8QoBqOwaQQLXKZYaQfX/Nf1l1Pg
OvdKAI/tUhFywJ0o5C1RujURmOeCSO41NO9XhRCGxbTLVMgcH7H5eGOS9nA1jgM2RsvzJ+f91vTT
Nij+WsBavTRTVqLUyV2FI3vYOwrP2WW90IbLZHYfSA7iYiL1zQjZr6L2455NT5c3clz3tiXOZnKt
3qgtTPTeDHzdZReKE+14iPG4L3f3KfoM+fRkvvnSWWMhpl4mEjLablDFWdBYNgwJorwjFwjWW/DQ
1Bbsufh8eI7tqPpxziwkCHsIw3ANlY153oZRQ/oprresvk+npumKsygqUIyZXWqaQwCjBPp6xPvm
olLelLrYXScq8Mz+RuOcdK03IAkiyYxMtP621m3k+3HXJ9RZZjT2F73tQMF384kEU9W9WnjK5YD7
9J9MCHv7VHpHq9jdgscwdt8ByNNS2qFrrtmt1Q44qSlx99rC17P6/IivqgTgvS3znx6tLoUvUELx
kOa2Oa19ZTIlPUWs7KuPx0UR9OVtAj8Y/k0WAuJJsc+fZlwUahQuKug5EyQgKb4Q8ayHFwJIps83
tgtrUafFhwLzUHSeiZjy83t2BdzvEF/L2rgkXvq0fFli4kmYIbF8NtqLmfwcTdQ/71BvU/jE/bDU
/QvVoCPjmUqmLZTMIfE34G2oxYWimSWMKCWWz2ogDxtwRzWjlsHVSLCmyYKlynrU9Fd16bpmTOCJ
UrcA3s2aixUVjFeqWlMSGXK1Ge5onQ3QHlu8DQLbXautdjPP6jEBcCMpszdT5dJ8oVv4shK8CV4E
joVHMvfpv9TGrlcVbG5OVNhUisF2CpNB5VRnMALnlakQ4s2njJJWzDCvBgje9Hb86v6w9hnr4MTt
BC7E0EYp2WL/ZQzf1uLqTzalqoaI//eNVeAxOcGYTvpa2L668lWx9P9+JogvoDaG/pOe9hpzD+Ty
AfuHn0J+YbmxgYM2VMFJact0pUDOx1ydclO6fQelO1/34GnlIQtba+OqR8sYuKgJW5uqOrnpL28f
a8I2uFebxylpdSUzkEl10uQDqmywMMHNxa2iqFGPn9Ujvw2uta71Hcf0s8yZuh16obbECx+0Kqqy
PTwvxIw1CNXy7dpExJ83v2M0Wlsd+ecBR1D8Ypa8N2qCGYKgd8u2obt63ysorIKCCX64E0sgkk/m
WUeNN7F5SrTWKbGs1KlQsx2Ww3rvOuD9l1niCerPPfgpS9j1EGw2X0WqD7IREOmEhiEaY8EWTxf3
tn5tRYAwtdHJ7vf8+7voPXSKY30EAhNTPMktZfrfElKYuhwEVBGAM49OuJHqjJeHLmGm7Dun6Jt5
EuPO4TWZsk4owz2QcIi5bAd5iLqB/A4rkVaOFXGlB+UFlOsAZUG+AagnLEwHDsNAaQQfMrq8tDhb
y/dhZzWaDOP3fDkgDntZEI8h5eCndf9lyAVyXjYieoyP213lrccFNqaLooMSNAGZApppTCYHeVo4
w+ds4QBi90wKZiBCzKt83MJGUAMrMSRu0zRrYZUyTmsXt/FRPg9mHBvHu7sltHQyANSkz4Viby2k
pUttwFGOC9+KkcIZ1qC6v6W1G3ZCmCqghq5a9PiivaFn7obRrekyF+lNcUyCCprSmP9bDDaS2KAj
6qSqGrmNcft/k+IKrB429gKhytuUCPc823556x38mW94DXXPukTNj07GSVZKv3rc3wcSE63cFd3y
wMa4uCDvWPUnJ/S/6xwA3zJ6d70cVnjdqJYAsP0KxkFLzwvRTnjKqdKcOZUtTq7QvAondXYX105M
mBoXOz/1O+MHmMLJ3u508A9xP8IHit7F0vMZWhSwW9wHiJWdbgmXz1DyxpGR9YcctXkVR/X2wDuc
Cc/K5gsTWjh9fSOIlLYMMqbE+3Q0eC90w8y3wWnU6ktMsRX/XohgnwnmaU/J1sgNiFBQMdl0TboC
QeyxmrNWlXvxRXKODCIWYsJuK6Q1/q6U9IC9vfE1Ai5/MqwtO/5H/JCQvPH6u+AceAXEbMT/pFfq
Zgylzy/kGCJoY+2d/fmGjiBSp1LalAmwa9TdXZUeov2kymm/lOh8/GL/mUGW91m15QudYqM7tnvt
3Z+AHN3Lb5F5BWd5GBenzGnzgXU1D80F6DjQLi9xfivpQ61H6iMWIFbjY0AfEQjRI8dbDIuD3Tn6
pigjiK17kUY/9wMga5B9miHGVqz0NWO9v1HCWk0hNs0QGdqP1MPi/dEhMYdkTTYrk3teWMW+DgGf
lW4cAWVZzjHMmZbJBnbFovZ4E2AVfvlW8OwBICckWz7qh+SfIUqRH6TJSIa9FFzdRUD1P4KBcJzB
/Z7qmsfKUBs50186Lw+ThEgeXey5rNHLI3Te7YZDvzQc9s9I/xekMqtFmllufdlXNE6D37eS8sQF
ZgVOC7Dk3xShS0kxUmRg9Lj57JtCp3z8IumbAfgysM/Ncoez5kGUKvg4Q9PIqUUBGnDj6XxzME2a
if70fYECNEZXCTteH0+Cjxfb/H64usn16vO3jfe+7FoMkN5MCQeLK6FJVLcqPScsarGZSXeh2Kqr
K3Qe+b3FmIub226wT9gSB1J0STjHVmY9jIJpdxQvnmJ3YcxC5PNTwnMCeEtbo68wmcqM+LHrKBXn
KiO9C3ypJNcShwiA971tHaQOl623QjrfHSSh5VE9bh6JfLaTy0k6e2lNdwvPP4UgbPo0U9JRR9t5
klADCYow4eoEzjcB+roMylTINLLmPYowqO/16JGhsPj86YwsRfkH5Xw0ojBgsrrY0Y47EABSCmVz
5nWWDJSs38BeDxEyeHhyoRDH+laX2m6MqQuAFEUsmcISOuY0q21veAW2gBmI6CFFmpLbmt5PiGez
n5il1rTF2At97EuK/a4QeayogzF+9lizdCN7JDUOxSDbIT2SBWknipxQpXuzzSft9iRTbixmzv10
yXwGOlbIfDGPiOuexcniPT0Wpq5CEuS2jfQyJwgwcf0s0qI+R+/Ca10a3nufg37V+g5JE3nl1PMl
eA1iy7PXeqzsog4EuK1jitOQsHJRcxKN8rt0LcYJwGtlwxgzG+qyS09ZQpCGqrS3A+1Ty7BuZqAh
0Pz4I12X/GG2znaGDzqE2J10+l+qQdGAO5hJvneD+NWy3+ezrXMpCONfsGoHQ9ufAPMwlrA2340r
5dBd1yrlqWEmbS8fz32ZO0705jMjl792WaudHVRKV9GwStXw5W5MrmoqWqJrQm7qxAeac2YQ01oz
JTMLfkWPFn+4yDHdcSDMpv/8npqGq4WYYhDeYm7cBZq0iJxGaXHq63JqO/v/6SZ325LA6IjzEiF4
SNAOerh5YiiabxIJPQFI5EJKe6etbtdq+gs3TtM08qTx2vaKxyl/ajk8lnIOu4E7j64i9QW32JHT
St25Kdm/Wx+TfSBlUvNhbR2oPM4pkqMqgVxdtSHunOdR6c1xHW+KFalr+Vdu1eP25oFrRJHTwouV
YLX/AMKVtkFk4YX2I/weyzhX+gV2kYR4gvRoqbAZis1YYlDK0AqDD4vII3t3V+PuPzTt0wYYzqG4
wknTOnDD2FKcDXWdH5eeMSzU6a4qK7SsZ2sqDHw6qi+nydEifiVvTHQpTpxw67FsEOwpaeICs3Wh
ScN8P2EzyP8Z7VRvPlrc1/ynaZH/+IPivtAiHKNw4gxECmGvyu75VbGJAaF+wXIaB/TqLcib8gX+
V9v8mhNYNG7TaIu2KJnE5oMHEEH2EkjwjbfpJHsO1zjOhP66vmcfpMR2SehRsynG8UdgdiB8loGx
ME/UlU0+cGrEne7W8uERTOYgbIQhZTbQeoNPJCmk3CHYxhtzZmrxV69/OrVU4KvsMk2vnUli+C3i
6W1ZAhN8A0h1R6ebYgEtTnGg3imz74HpSh3zZJA1kCc+pZLsRW7wsMbQBq1IG98BRCPmPZ8Lt/FQ
a1y3GzRiwC3v+o47nofH21V+UZNvVl7in2nJFDP7LxDFlaRq495KjC7h3skVWi5TXp5qlyfUydU3
oQa0DS1wAq4hv3lTOeKTi6oHTyC/vGKC+0E7HY/uGf/qFAkOaYQ24jbHxNfBTLjE300VW4+F6R0x
Utfl/kLUX65NsZIcWmsLUilKH29ehHE2KwWshMpWOFDFSBlnQaF98vPJp703k+1IL7tvC7p44Iwv
ou5PAH3GVbwVDZQqoeGEkRts4MV0VdGJ2LkkRwFFdnQ1GRT34Il+k5EwA0GngkZuFzXIlofo1Qax
/jEerirP/BFhxePd2IFfAm8+HCXVo2b648LgOcwLTJWV9WJvlz5nhpI8Zi185m+8d8WTB2rhzZNY
xNTa9ZF5wiCntCz1Sw3YOq/lTWEUDANc2rJBZrimaUwHAhlgL370V125LRac1SV2tSVBxI3XtUSa
h+Mzk7T4raW8TydAElBiH4o2C7PRIhFArs3mrONhpPI9zQwdjH4jAv9iqrEya/ZaHgXhMba0XnWi
Kfb9jhjkugPmjA9ynaKWMm7dpcvJDF7TTDqJTaaHOfu/VTbfKH8vdweNkN8LYnSHxKV4nUtLqfdo
VxeMUfBYnP/c7ngXKnmqVD/CBl4th0bmZ8bV8QryV1USNTYUgTiXANws/zc6jiQ0rBK64NQu89ST
ZN3uPJfkbVlKfvvat17VXguBJ/QptvOwwto4bDRTbC6Uxh/L1R+M5kbUERhnIDmT23/louuv4qTK
XQKfJiw2CQGpO4zJ1bonNJMbxXCclhOLs73dqJLYEWANdU7TfBadncCJm8o077HN4LfuvGELUeNE
8VL54bHh5lIA4ghlT5F2seNI5NoBpHTO603uYkFz+oTcTbOzvfKqBeUfyNYB7OQXXHYKqMojknyE
v/iI6CcFXLCek94iD9Pj4s6zvX7twXfTiJENJkzqtGegp4vVjd744e3zCwBhChu96vin86zHISeX
TaGQxD+n0dsnNXTtDZ3A8t6yppsXDoqnUAIXX7GHUDuwhy0nbvFx5iHZlzO95Y+iDR/z3VA9oFt2
+hbliWMLg46xYWkAp9JW8YTUidyG60fUzRHnFU0dtqmofGYxIqMVDIm1i01wSxZXeG0qriAAhQCM
FD/9EBTOR5WaLEZTuOoffnK664kZX+g9/fIa5kHvYh10+Fg8rmDVFn/Z9/g8IMHc+ds7xprZDzJn
e+mhLetSfsy0MCASnwsE55o4S0XOBBd7GIdy/EJe0T/q3JbC2zgq7YHRAqz4LjywNtRnby+bLZxO
r/5t2sXM+oDv1pRsCDhFQnuCRxSO4LuXROeiDUehILz3UMGPSvGvpfRfyyuMBnkjqgm5JiB+H1gA
8orzqvKNvpxWuo6BLgCuxfjokG/N412kFlnfKWBlDwz49oQnkLoFr9sUaa1bLgQIATFKqFsKEJU1
6tNEHtlcmEfDH57Cmu5HiLd8ORU30F9XJ0wZovGzgw0z8syt+olc/7F9sGQxbjx6fmXpu+176uTE
BtunpJAsbdWvri9Y+XS52GPNAlvWJORj47LppW/dMhlIE7mI7z33Ot0OlnBfjKaBWHYkY0WXzu1f
7l77Htkz6TXrcc1XgBJmGuVrLstXAXICc2qB+bnh5w/7O1Sk8jfwZ18V+1VWqEW9fFFPxCzGSUaM
A9WAu51x0OfQurmQI7KaB8GGmP786eyIV0iN47a1XjIuez6ilipcVNes//7SLX48XS0f5rqT49U4
Jt7aO20XQ/ETGOyrMcg6SBI6/kbHvgjgrNotNZ8FPWFT9EmxG/FpE5qkj3mNvoFGa2zg5N5gt7o+
Igp+yiiNS1IcfUuRjqfP23ZCdpF/KgHG5qpZY//Cb2EAkIE0nv/Izm/R13LB6q5eXwbv/SGLtdnx
To8lNPFFyCg18pa9Ba5LFHoQ1UceLswdFcoSpnDHGUyXe3E5AJsGEeJbdrT1M6wlAPknhyp5LzzC
Vs5BubJO1lwkXlrO8zzJIItB2JHeJGSI+eTPialWT+Z0lhvI9vYURFKGiCpPcfWQ5o8EFgRnb9Bl
g5sLgHZ8d862SqYx+mw50X/2YvLOSzR4cTlZzayifhon0BwDb2Y/Nc6IMhPWgiUPK/h73b03BfMG
7c1+pBc9DbbOv9Pf6Mk41p4r9BciIc+Gkm3myu08i2K7ueU89EUmOutIb1IBRwO3xxXg4MEaWlSr
QnpJghCeEq/ok1+X2fFUbHgWpkrLuzYW89EUjBzVtO0bMdHc7cI19QsRvzkaCi+9fY8dKNnuot8h
j+mjGFNcuzBUN6FFsP0nUoOH5Ws1AWvdh0/KJkh3Ma/XGpcwoBg3dTVuWwGyGu8fhedroL7teY2h
dBeAPw3sqq7lHudlBRihHZuJNZDPM7mFUlZdNA4t42UL5yfqShTTCaw7lxs1YiRo3C2hSwLv9Yg7
tq6c7pfha9mzg8/M4lGPMuyKp7qfi2J3N1qNAG+nl9PZ1tcCX7WQ3AYif3cMr1j58NX/6EyaddNH
4Op9nm+SVJJBy+fFOL1TVUAfIQEfZ/vVBhyViHoKKPo6pL29rjsjEaIfuN3ThNvMLUHRDYqAHxdH
BHxW2miolZxejmObLGIf9s2hkRfwHDXMHot9tbu4yG+Xipubh8GiKe8dCuVb0PyGls6BSRnF5m69
3yQLmtC/UF34L0yHOGAjfFaVTzBeDjKofcsusO+D9Db5iQkpqo4tQGiwwR/4Ri9Awyi3+SDJhhz6
MEij3olIbaZZ6Z/UX0OI0jLtck2+J+wbJUeTaan+h/cZCi9NTUNnNxSZ/SZHrd7pK5Q6MKSsXPLI
my6ALYOL0GvUoWt0RHCIIuYzxIgKzwXFBP7cbPZ5LmINWZVphGX23CPqj3Ia9TXp1iYcW5utKJBU
FNUIedAjJ26ZTeupML+y8JJztgKdhOrd67POz0H4iPjVbdb0zNjhSTITF/AdYEjw/SSt9TBVp0EZ
w9SqZHLu+Zj+WWEJQ/kIaDMTd7us14QPy1XhsDBqUAihPTVvbytKju2FqcmRy2v1BAWsocxEc0lh
J4i1Rxn0usFGQ585zDm8GLMoZzvqgF0mGvdljXe9UdLKNsZgSIFL6v1CRt7hETf+DQdeqfTTZOcI
g2z0hs3nOJ6vGTAIgp94sXNL+RM7KOPuewUAPjHN6djImJFA/fIGnBlu+Y785ClKK0y92ycVCdw7
lDlV9o/wktqa9dkfC9KzDwzl1VG6BIwU2q6DY9ADH3U+Rgx7fCkHJJw0rr5/ATqdLzUpsToz2R6u
kXqwFWZW53n8HjzWxRvIEDy0EzhAHgt6V+ODvlt6KNo9lDonY5nBP2MleHhevFXZ5H1Of4YX8Za+
ERJzfn00jo64JZn7XZkGur4ZT2dyIKztFwaX4r69nXcLBEmubW+rdQUX1YFArUF+DOFTarjaXgrl
TZHwegqklJBOXRmQ6fFxGx8OyF5OZ8sKsHLw8sQEnTfJMPDRqquC66nkiN7Nryk2uj7wkbLxbBEi
AXsMJQfA735aWzC9uTL2s4mU9QBYEixcFAIWBoI2cbgBL8TsdViDJcNt5mKP7reMeDyHNDxgDD2t
o6mrrpS+glLwSJHYtDAbEJs5tP3Bt9Pa1l+RKY9xuO/pHhZhz8rB72hbS6CumyBv3o/AtuGXkHmX
Y+rQLGJjrib/wmlB0AcFAI7aAw+pAVow1fpSFIPXo4fDIzoixoZtFHAA1LsdmZ6Mcin+tryQ1B0u
kltmfZwqbocNV1B5cakg3DirvfTdjruHSxhy7Pis560KGEP+YxzZ6FsDP8iWoXyuHNbUoXIpWeN3
MBsW3wfd9F6G6ezDW8ag9k0URYCuWiqPUSjjsTcVMcE7NHbD1fX7eqClPro3DAKwhZ4Ajzo2tqPi
VHig59D3IwwJFMhuYPzSKqmJhkkYEOyBuqa6Tvyb4CMiJSg+A0bcU6FnJ8Bqa3+ZTzgJjIxjrFch
3VWovrBDx1EhQQrkQusd3YnZIVnBhcIUSNSIaDUEjoAoNLW975Mv3mi5ABadwX50CS8SqxuG5svR
YoVPJDOFJLFWvRo4AFd70vW/U9uXxykG3oYKn2E4ZfCVadmVnBs0bRksbtphlhkpVg6+aYIvd8pt
39TfHlV4YV7cfc07S6kwhWx3MgwmjjcLDTSGsIjel6PIp4bVH6r9K7I/BIAB5g7xX+6MGVtJQ6fs
ZpOgZGgARiaw6uUHe0yGoBSOl2+EDfBLvio3+ruGwV/eAEaNv3FK/0fMnG6apqUU5ltb2fBy/RA/
J8JhfkUAyNu82hYXeaW2iLECZwYpfU9ZLxtB1aLIKdobCB4WTjZrRvRu8AqjYJgcKKrfbQY8tb1H
he96ZJcvVL0PzbiM7aM7cbbROoVQNvWVpDV8MU1HHR/5DqAWmTr/Z8LUYzuFbycKTNUpfM+p2JgY
xP843bjH7wFqiXT3RXwTd2aeF46UTZmDvl6qML0nwwzdjwGV6W2Ydjh3xk/zSmNiqf1PXseKWl4N
vQakjdgtXyv5cJIulul3+xOYuaC759UITu9Gfm0ZczOzTXfqNPMn75vFUnCxepKf1wVm4y6rofQ4
rlpydSnFp6g3nbKi2s5rvw0EHruSM4udfrW7+2vjDO4spZ8zFF7O/GxjcJtamURi8TzRj3gH4tBX
1JodOizJ68vJHGNdoqBXFhF512SZ0HpEDgLEuAXJzLMeBag5UWD/ee7S+K3MRsyl2L5fpIf5Hf93
npJG255KVq0cpmvvxgSb0V3sp/tQVrLQ9ziOFRoSZio9RlCSy5n1fxMxclnErUL5sMMTVO48yzEJ
PQgd5XBPJFfkQ/G9FJc+uszTLQOmfdrgcfJEqrft2O4KucohgU9x+r0E7jjJFWG7I2AWvwpjxu7F
QrSyQZF/d4jSwHMTEZliSEDOs4LBo42d0QhSW2joju7fs99LggB0CIxjYL5ctAazqoMxlGDyjVxZ
zsaQpSc19fbWkjNAapnOStpbOLlacFqS4jW/m7Orh5AdRYklaeMcLq/5fTfLCCRBievvXxhDNy26
lM2EzEZMQKbddL6tTsbiRvSQbprVdx+LTrgqVdLe54ESLOdkAwppXtm27CPvfP3Q3ItUgPFAo9+k
wo675RFidbtyRqAtO7s682peZz9H/nIyyVj6ZJmKpH+6xiWKhAhSA3PZgU6lYBQF+EN/t/JXfPwu
cFDP8F69SVV6SlbtYMkyVcrlly1GWBIPHmBDMM/EhyVJE/nGlYL5KEItKpf/2XQCc+L0znez38+t
rID3j/tXgRw43SosHNBaFSyVF9MQVnKJRPTpQi848taombBx9shDH3illDukfolzP6Mr3Fb9r8IT
cK34XkL5ndNgoI0vrZN4E97kKwIjNEm3rIx7q1TTqY1WEArNKgNoir5bUZkPJTFgaFUlT9t0b5mf
Z3f1WlKVtOZ0uXReZ5OconHNoAt1Su254wQPcG+uygrBQS/5QuQJmTrDpM6llC3os/F2U0ZTqnmh
6g7OVaBXfNZbpmar5XB79e5C59VkwKW72/Zt/iWHUAtecNtffhZotMA95cHI+0d8WjdLBAuPiips
QXiAVOCbo/O7+zTdDhMYgzazm9ayJEbf0gm33lVc9zdjzqwk9WjnPlV8Sc6vI1F1MbllgnoqQuC1
fRQnqN8STyYnpgsvkCpwjSjmgJUT8yHVR8hWWt7RUTeK/9U1P0FYQ7eg/KR/bHfT96qMniQ5BmHM
fYibDGRSapR3qoPHIy7Go/xsOMkDjEhNykwiQFv9BP8jhmSxJBOPYprNv/2xRKIyYYMWqSlNAfiv
WbypsJWwbsg9xTWUVyEDsrv86b5VR1+ZgDmUseW3rtZsYDJAiBi9S3ax0bKgO2Yp/5RcXe8os7Kb
JjpZaXhd7uRNK3bt5pOyWmyl5jPpzmS2OIEgAvuxsEQijLmwUDkhx/qH4Haz3Te/jJYJa7aAGldv
CfaCJgU4654CkqIhBSr/GIl/vm9WFgCjWQvO4cqdEp2xlXE7Z0fDexKi9kz6aNbAFvle4ZrWxPkx
qk8qGSKEFpKvOIKm+QQ/WhY3eeJMui5bOtNG7suMGV3ytm7lip4N2fsWaPrJOQ+rxwoXW/c3EtSj
LeGPW0sI5j324KJ3vbAiytNG6VtIULDwudSvktB6VXfGX9RGFeA2WHwu4+2Qk4NJ6cYZnn5Po32t
6KWsAhYThOJELpcYwO974XR8D7uUE1TbgCeWcYs2MeCt4KsdcTySHZRkJ8dG9GtpWGVk1H12nWRP
/WEeF4nvA8EU4VGXAdPc8611seSBIAmOgr2H88igHhkyjLvQEVcYGC96SODrNrDDGjyYfO+3H6uE
sg0Q/V59VdyWyw9EQNFKtPZR+3MMyqR07okl92nn/pp2b7PZPZ9sSWcmY/7MmWKQ5G+v39sh+mgZ
2CJNBxPSnUxx1fx6KElqOqWUg64WtPgJBX5nazpZ29xzDFmg95praGTMAHanURMSg0dXubAf08WJ
rxjzXcK7CjZ53z3jwtQ8pNnIph5HoLQ1j7Jq3Ao9aRItThU0gFXu9Q6i4vIFVzkPZwrVSonNOx6W
5bJ4O7/LxSTJqjoBRpFRHkr3VwLZX2BUf4o7gmnNG2pE2VcJ9j6uj3iNwNi+HJyALxsswSwVOlQ+
xl/EkDb+Um/GFJYFAbT3OXDVsUeawDajwcajyF3U/p+hUNbwQhkOdIaXrgg7HLm4St2IdaAZwL4j
Gq7ExzprR01cx4/CzP0dCZz6vjWyL329c2dbFaetx85ch//BVmmuTiv1cXKary6BzWYXgHemF5IY
DgvDKytMqBwnYI+ah3JJ4K9bQCEH6xAjhQegnsiNMpz6muZqai5w6ylsu7H0PXNFvjGKo/2GFqm5
cCxIVpIFvZGYXKqLJWoqEysDJOlu2JS4w7R2hb5ww5PDB9hnJTq06UZSyfQzGtAmbpH774BaTA4f
IegGZhaV3mkpdVwgxE/qBOnp9jnUNxdsFohCxxy/VZ2h6vGMuKRty3K8j00SS0/KU2oEZ7na1U9z
Gnu7Pa287LyA9vVBPLiAKtYgMCQGZUXCkNqr9ABXP7Mk5RXmBtM+qCSqNS/9+RLx7aWC1B5F1NtF
/qEVrW8My8JsubSts8WEj2QWJ9k3POL8E8xsX2emLNDB5YfTu/+QHMM2fhWcejrp0e2UO8NoyN3Q
e0Kri6421W9wBtMJD0mt/JIxVrmefHJPlC8nrtDAj2nGjqqJtluwIVf/STOld0qabHueIAyseKis
kO5uNQYEVNitm0NF5RKC8zIys5m0tQ03vFNLk3DvmT7h0WvTJ3XRia7o0jOnkil+49+qVqKmiI34
FK4YUH83iOwc8Dhs8I/2DkHXAikaAWkG5lbsoRrwrkoxFjUYY1oTE8COhEcwbeDxWZ8JmagyMoTk
ldXMj+OSKfycPk/YdYyQnVIN/juEYC/2HjnU+DC2fwik/oaDJllv+niRbsR8EdjtehGIaxz5kj64
/Y79U2/jvMd9YQoCDtbETyprr8ENMDHSW0vOUScfVlQaO2cfYaXCJhhi5Z0cpW8tlAX2izR7XS0p
lcVXipMFvwGMoEWn749woW+kef55IJBgmoOeEir8CtDqNFMa/WNYjZSRCry+IPhdfrf2lghV+8p0
ILwz40lUpG8b7AsFz1DJSJCf+liTKd2Tn/wAtdk/OZ1abCQTzD/2/DloiWy2ca8ICJYBes6/ZvCq
rFjwA9tyQiftDW7osKFbJyqZzAKP8cJQ3nNRJPga5BDTKjpO1OreiD9/9KVbQamPITb2FQKclVKQ
qBGlPLkXLQJG3j83FUX9FslaCQ9SUukqDJDeTd+wwjWLiIRamj5KKcIJjdNnWMbf6WVo1gmxJibQ
dADDcX4dkVwGAjX25Vq/AYUYomZ/OT00sA75wodYq9KNrhl4a8BE4x3NQnZu7fECmC9wICDAjY6Y
mwHXhhRZ1d+VdA2lamRAPuPNiPLKKLvmRKIKUiK0Kg9OrnJPBXLCa2lXcbRr5HnV3/NkyKCErGe5
S/yAsNTXT98RnxhzYHWAz0GRrBwyprYCW0qlGXI0gpBsh8I4JjS4yotVYWhCS2aHwIGMUk162cat
Dbic11HpmgVTiK2LTSc52N/XcEfP/ZYIGZf1nRXQuxgczu1upD+0FtD3LLebNb8z0SFuiNg4Ubkm
h4WRL+DgGedTRDEWHqpcFsCGQe9dLI9fBChVSBy9EO3F5uNbsrHj9G5OivoBUcAOpzLBmUzll96x
pFts0EBMM3O8ZpHETpc39yu3/ErCMiMbY645rLdX/GdKuco9r1bRDlFkxuSrOcItTp+v8ULbhqeM
JPJXFGnuSpnj/BuW1NGBpIHyGuo4HLKB+0lT4sgh6PjJrxaO3idM8S31MNjoJqY7r7dICV4A+/x+
GEFoyHdPxFWiHF7XC4XcpoQCay+b6nIN38mgBn3n/04i1JkxjKEqB0n0CeLqi9DiTKUsYtfJgXC2
0j56RDBMY7r9rL8SEC0sJKJPKZ47anJSVeOm6AeL9CyYw2d40l9EIRYjBI8ZvFwQ5o6ZXL+EpKKv
grp8pBR/U8lTN1jvM7fhwtrviJZ9W/D5qJFYtw1y+ej0fFhZLc15QbzBzJTNoqTkT73WWuLBuzOF
HzLdb42TSL41/nglNX8J/TpTsT2rAgnelXrybblhxP8aCAgaObOOAuYjl2qrNR6tYtAM/0zfcIet
5j+BaEjRglXeSilA49ihUGhgKUQZcOSo9CnJUScO7ldSSQiFMd/LOcP4C9bDvBfv1ZEB7Ss+os/e
ZtuYs/059t3NpBPWRrog/03eXhaeHYpw2NPaouN2ilzYU1NBcGrV7XUlwkxlQvxOBLegUCsA1a0v
pbFqK3G9k7zqxflvQN0EgDqDzDjJcMGaPVdDgK7BkfFNwgeaL56rW8jNyVCd4bNkQkaMYterVmnX
0DTt7VFc2U+Iqd4wt5sLY7v1QtK1SADLnFGRnZNusF1z8ny0ZwjCwDCpc9T292B3Ie5Sm7K8FVCz
/9kTbdVhShvxcpLkEpqxnPsezKUs+cB3plZAHyn+28T1gOuzjwtq6xU/XUGzQs9jaHM9L4LTBNbC
64s84UWUdznu5GnQWqcJYM4m7zXMEA29iXcPa5qWmebGj3La6PwxlhsBBrCZVoiV8lSKqoBbtfZ/
49MtByT9E/LnMqXbLJHfizifi9iyPWaEJQxmQIH3kKwrMuiVXJG1CZY+54i3yFfxH91f/aXss2+C
OVgOQC5KhWSqgeLzomYJ+VtwJL8YQysa4HJnd/dmB4RbBUyF8Z8PAjVL4A0mOBdhN2xMoDMqnu59
tZK6XvXbA+PazqMpMyLA6C+EXLSmwOu5qMm6qR39yV5kDcn2BbvBENNTBQ9U0W/ZNYmWY2toUiB6
Zh9UwhbUKjRDc6LwsheR1o991EZ9m+7GGBDCTqjkmj44WHetzmuJl3qGMQXgI3CRCeU87Z6Oynyg
vpKoZZI6/uFRXjfU6yp1XKvIs20jkjJKpDv5gbTDG9itwaZzHrl+pJw5tWulDPtUZg/nk0vu5qlq
NGAukNLjHblg2L8vsP0FBBwIM9c14xWb8nZawBywW4dSo4lPSgV2f/e4Yr730iQYxzMrkUorEMY/
MplaMuZ+sKwI4xuXgVZC+yWxGk3CH8CibZcIuf7JC5r722Sq8r2MRgJLKtRY/GaXtQXnEZzGMCTV
cxrAi50Wl6IV01ffPDbzn4kby9IiXGp5u6VdeydTmfsf5UqXz6DprPdJypARYQJT8E0OG9aFxFP/
Vt9KxQPgzCChAG9oaPTXnszC8EiqgDRlW2CyvCS5JuyYWXHiIxerd4I1Ni5bNLm2BYHmxvY2ij0N
ObSaoXFGBbfsUufZQxDLk+bbPLP3m7tokPJabuk+maQP3uz8SFgKHIkj1grGWc6ZibOIm26h7oZR
g7WKEnhEdfbA1OVaglpERuEUp8ytUKAgodIPX0JWTVqw0wn/U0HFgFteT8Hwwll0ol50uDYv2SRV
eYtS5o1AmPK9k15M5cUelAE67rWXh/uzfJPcKh6Th+FmdSMbx0N6HvMoLXc5sSSg/z2Yy65itDb1
+CF+5d0wUxGXUywsecgluzMq6F+jXYcUOT+BDjAQJ6bOYQ8mUUCxAREUrfRtENxHGuINappa0TT6
uBD9rYvqNEJbelKERxIJZoPTtnCszWMLkuhqKdeLjwRS8o7nBm7ScElvtipn0M8/zVYyuHJht/et
cf5ARDlhoafba3PmXUSx7yfiY3pj4V8L0GY7NsHedixKK8W/2rRzDhQR4ymSmxu6y157Qu9gns8C
B17kZALXow4BtmpC5NjgK1XiGwN/UrytkySmBK2FQAnNgKqIB5Jo6Vph2bP68OpVDT5BaGHdkTSd
HD8rGYIh7MkBd0Sz+n4kCr1iDiA3bm/xF1ia79R4ptkoTIq5eWgrTUzvpKxiO9J/L/Y5k/EsH/et
Xc6rWcW8clLOtuk1hG1jjzQsxeRgqlIYkvuUq+1rem/tFgDPjW02QCE6nkvA1lr6/Lyhs/hK2QVg
pAHzCdoL3kQWNmGOIcsGpBvEJ5BdrueVq4425mLlbq7x2lh+Fcx4Snd2eYJiAsyx8w4O49i+YBGc
o1K3BXIFIkQk06Vnei8sqwEl8bp/WdQCsrJSXi60uazu73FckAFb9k9INSSI+L0TUmWLRAAIdAAv
O1oGYQssqGDKr95DGSTHbRfTDBSw8M3RLefG7P3l5hidlXa7nDi1gY0aQ95yzohhHTO58nmDog4K
nEz7PIJHZAeF8tLnJWMg7WWYYcRJK0uzy24vqSMc99BeQEofUFfSRdpYZkoH081/1YkLz5Kum9jc
Vaav8V9m5kffc8S9WCFpNKvn52JB/by/tYo0zyA+yb1IsMXW5W+crNwrYuop421np7xI6FSzJwlH
MupDiPb5Mrg5kcyN7BlKt9ghqkjFA9QU52yjpLgPNBCfsYesYsDxK4wdJd7Rgs9EsH2pl5CYwtAJ
+LWh2n5U36B8YzfXGCqxhhx3EtgybVpgDK/89Zd6kLvjpLCGWYroJr+1OJMrvwAgJju7S6BHtx9w
7JUABIoIWW7zFeUzUhlSK1KrYsYqlADcq5J6b+rITknSmAKkyOWR84nPQYkvbCYAMWNN6gFoMmc8
MErlhnw/484qWerZEVLBR32kyWsh9swlOxQIsSiYjGY4jdEUOBmKXTwfWi3vd1HT21gqhdFj5EOy
BO6gGW1JGvu+0aJS7nERuWS89zWZka5sh/eXGmL4Q6L4p6M1+T0pWWOFxXyas2Vwce0GfBEZfTSY
BKR8h5LSg9+l3Cw4bcKo6D/X0TwT/1OyUBwe6ceDJwGHLoeHoDaNy+Gx7Cy2KjK82SW+zvsloaPW
1G1ngMlkxL1JHW08SBz89gHN57gozp/J4XxgZMJ5Sf24MytWZbfqFGo7d070ucck7j0J2OY4f+d6
ENt3qv+K1WlIeA866WALVz4kqFEZmsCPmhXcziVHjrNi6N6NVbjagR5uiL7q1UHVjci/r5ey6CoT
jaoICxJ+hXa90bO8UXEKgT3B+orRBut01Xxk9auzCyHN75PwZuLdW3gSR4DXD0E5WD3ZHR77tsHi
KoU0VDf88KNKid0jXFPxmMGW/iPh+ijxVuYt21gO+G6Cmz6wrm7gQYNYcnyrtEDEmSxdv3eplVPc
2hiZTQ3srMwHR3KHr9dWISUkbvEP+W1SZfffm/AA/LUi28FBYbkRgDkyMXZhenxqjiRYNzWutIST
d83m03lAxW72a3mxp+WuTkam5oP4/Im17mnXNf3oZxxmm/mzwNyDXAyx9oOySP7ueovtxTsq/z0o
bSRreH2CgXW6PyhCZpAzV6Iq3syA0YuvvORGdJPGGo1XAauNe24gtaPNv2/hrMnd/lXYHHlbji+U
TGJxApd7bSx966AoKq+Ga/S0eZG8RxB9UpnDk8bUkXPC+OTKr50OCXuU0kVb4HRU+N7TSeWLH/F9
5AW6umqZszqdVATZq60+2A6FKGX9QoOr1Tlh9WkWu+9W8NopEMwqzAPx+ENpIOQtU2Gz7erBooGQ
SS4hXbdR1Ush39hYghSVw78PETu+0Sa5vW0gWo8s/VGiwSBQt1WICf3WpI0DMalajWwuy1e1AwEP
hwrj34wdb2R9k4OciJrv4z8odqki9s2dQ50aPYz7Ilx0j5V8LN0UaRjuwyFGSnDN1rFzhvhMP8VG
xGNCw4i47KhG0Lf2cZ6OGv3NtALCHxxyyldoss123NgIi+0vJi8gfFxiQWwBOmjms7FFByjVrqBb
9tf/YHEyDsDG7c1Q5GbbUDFJ6ER7t2UkvYjpD+92MsVDFrX57dMOGrOLPPduQ5fYTWg4yCu5KM01
rE/XhekSIpyLZOlhOBOx2xHm8BmAjDb/09QzuzbYZgQGRs6ZGxdU2vrPFrlRAp8j2VIpaJufwuQU
5cea6jsmqPAbWnXOCeycTtJ53fMaf4u8qANYxa7NPngG1r8z1HzmBrnPazOA5EIyze2PTyPv9s5V
bXWGH7GMr25hmNyUrwBzV4rSsnrXMyQn0p2d1hZuYNsbrNfWSLIpLYfFu7+QmA60RuAwxcFdI5of
iYQfUKUh4enii/d4XZCmDV1/Jt5MT8chRAT41RfQ1EDVrT3giCohbmETSDoDL8RldV5J2u71iGcN
2i3uQUs/dxjH77aJfPT7RwjH9/AO3RPdWALU05EzYgrrNYXmJn17xBp9gPXKSObOb2JCuQKpWstm
mmlV3HIn2HrSPYBKZav3e1RjW0WrFFXmG9Qkq1thc3wlQy1BYrgS65lHrVPQ2Jy9AsTnd+JHI8Mx
jv6zcOm7FTpDMMjlQP4oWffsw8avgsCuT4/AmtyPJuMOa6Q3XXBHc3byOkFaCOxvBVQnneGg+u7Z
esQ8Oo5b2OtaQ3blEcHfUB6dV+4Ex+kZ82Vxw7kSJtH/sYlkYHiRKYsNlyqAISmkYdwJWPgnePJS
7TvBib7s3mCU8qEvXkEa3W00V60cR9Q0VrXpRmUyLFW+q0C4GeNyIWZB3Vx0URd0iZb6SY+DgenI
n7Gl/jkPcHmc0fszdXk+0VLsPGPJixZrUwHJ9xJuWiodEjAUYofu9CWYFh2SwbjSQKm1YicQVup3
23QXo7Kg62kk191uGoilz+0+zkQ1q+PJ+0mAfT+9gjb06wgULAdO004AbCkbwWkkhJO4tSiE5mFO
xr99fzuBfWGpkX6zlBf6kHCp5brY/NXHrBl5usOCqZmp1MdBITLcLN8p9qG7jvgHDlX5TY3i0WBr
CZ8/qN79cMEOEB3PPc6XYe7oIFbLjIj4zjYxGq/MmUKScTuI5TPCfxru1Qhu4580/7kyKW2eOUuA
I8uQqTBfgNyMXYxsIyzqLC8B/8sU1INVaWb5i1VW/nNMDTJFf1P3PT+gv2ytMriMF7CQyXUyxF/q
MKOPnlyL5uQH1ADckCJLkxXALBYl+EG7agN0R4nqxOxFHS4NeU81u5Vt5m4XqKqiRO/nwq0LHyoz
r1sukwc2ESEbKpGj9k8zht71hfZDKhxlmnlc3jGXd7Y+2I+mIMsVf00WlAi1V2VZ/0OINnosyVlm
7jqSpHRC/QK+PcuEo/4D0PEy1M5Nf6eryAnLkV2u6xSp/H8V4+9nUVB113CUWGRqjnp5+vrSaACg
DdC03lU5MF/I5/S0D6gr/YDi9FrouE78bj23nQe34yFT8fENJTDjo56Ip6Mbaa11Ifh3HpX3Ef7H
xd97GTl9TmQwWIXL+omqUjeS9XyNRN+y2FnORumCa9UIhQw22vNsK6VXwZ4iZHwnJRK7yB2npR6i
G34AUFzubCMgWxot+gkkpZAzcnzg/KNFGfRM3Vg6Glb2WJh6XuXk7GjNBulMlRNbRs6Ayrj0L8+a
FdLBd3Gkp7gm4sOR2qbkgV7Gqp27sxgxuBlme/Umu30det0E0le+jYv0AkqVzQnPmAuRxd48kxpU
vZwI+MkC6lPJAV3nPp3ZbEtJrTKA0u5o4rTUMFEX+/R3Zn7qOw5sFSaw1o+icC7IFLVKKFm7on+K
u0ebR+SLVTD+lstRvDkjLVqQiAQUvdtq4ZJXFJh0j3rcJ+fc8tXTHf0cwW6LyM2fDs1u8C09b7to
WDTaLPnEDKesjafSiHfX2tUKiqKuZsW4JN/YuszMBN7KFqm/yJrp85SCeV3rwEqmTwhKf4IQB+K/
Ht/g20Ga503PCFBFxnzES04ks0P7o35AkxhOpkvuP9LpnamrixYEqCIAVtyhFFDt3Sm/pME9LtS7
9Crp7e4WbD1qrIUrAmzLWFUhfZN4Dg6T0cTei4Y+HyUdS53OzVwCp/HOQ934zk6WES1h+whGrNLU
LldTW1KTbnrSNgvCPHV/ww/XVbomHxCgk4qH4bOhE4eSKRF3INxIpzzz7ZLJKy4vmbFOfj4LbWzX
9XqpnIKrHye0Y7Q+8SyzkO6L5yvous0o5YEXL5EaV7Re5M7ORAS1ZVYuNpsOJ1qbpUHUcaYpQwmq
Coj2eKkLPrgIYDGe+PwK+SHZq94Dsigdg8P7UsGxiMeRqrepal5Xe2fv9MfvdMeID56f3PQVUSya
/zSu0wY+7dMI2lqWxKw22yseVSpf1sXadTuKjMEp4gorgPPThpVA8D+aoAThzulMQVaHQZdds3ga
hIgjFO2WoOptPW1YLr0r1iiPV3eQyShm1Kqy20FrWgpMG+fs3lq2+bHeCUhIN8ULQiDdWY8Wge+k
qXuHp2Wzj9fPvFAWiYAlCGPP7Q2tEO5JwehMOgkfbHJZTH2tNhEzzxGABYl00zs3w8NmTKN9tyQO
aG+rTeabdX7vtD3dCwhqPYh0+q+LtYOiynP+TGddIOc3M0W9PwOean90PYhILWP6hbLa0w4kOloc
+YyW26dTZxEQk8hwRN1WDTNaz3WhVXx9rveLeHOQ7By6ZVTmQZngQXQ/c/W5odqBxVhlPyMMY0nm
o4D6EXKaSF89mLYiqqCt5L3fqGdTktsrMw3vPQIXgetBMJ/4j+0ztMQdhlMrL/+UfxiYH1WDetMi
WSwCPrdm1V7gnTjn8PSy327c/ArT9vyHtS7O6LY2LVdf5W45ASDQbBTLrglbZNWBZNOZY7lFh+gr
cZ/XRAO+8mXzFYQYQAVB70EQMjGl/Gax4Z7ohrJtffBC27jw9v7V2XzxyIQuIhjyvfNfYU94C+d7
+TpEaxf4X+oXYWf0egzZKQETf4OVbqeuNzM2wJXJA1Nt2MlWAZ/ATuW/eu29ReVR7pp0EAI62JnZ
hNKt9cOMjABC8VL4rrINI51vScLGnhySlWmGfyAgSfcCnR/YxvhM6FgaPdg8oWr5goL/sSdQQqqX
TJajVNGnMKn+ZNv8jkY8ajTrWoYwjxewOXg5cGLhgYVZF9uz1OERLuUPAB2ZIuvBcEXsv8LRApyk
yUKRrVRlE/lT+4PFrPIYm31l9N+gLnC0t/AwAyMOWpc1yV4cna6WxyDYT/4D6E9gncDJab//eszu
J1MRa5qYiZx/HDSZc85OlDyXYHU2NTeZ97sPHM3wVMnFl7CNYOMOmd6sTJGiuGRbkClYz6lbRO2Z
g8MtFqu/1e7r1JEY8t+GungZsH2JmVgb8VshW2y51bHy8AWC00oDxyM6ZTYOlZEzy+7MPnYrG7b2
HXdJFXCi71f3pXR1EcPPev6W32SlUNloTui+/m68eevPHmuPVUbyGfVKv0atZaRLEjblAobXYvZ5
USiyBedOCN7ODMNRYemYHjYQ7Z+8IZTmClFyOG3SAmiWUVfneq/Z5eY3f5zODYudvgw24yF+65ux
KwQguE9IY5AEiy6eE5aBFlh3VlxeTjNa9OU0PMvIUO8oTr0qP6QhaUZ6rfS2yucWmB9lDQRzgvgc
Wqd33Ier+elEXfFx1ppq2YCbPGz8QBESE99PniDyRqD/7rtRSifdIBCzB/5QgQXejPNeA5Mxy15H
ugEkH/JEFm2iviuVdHmI1w2FrKnDV/c0jaIk6b4xvNIPpXcTs3OAa3VTz6+tW8CV+SMUsh0RcBAm
ObUf+Dh8fE8QJ9EterdUFfM6/A70o+mp7+FAPgxFgbFjXgI9vDYVrfMiCxY1v6uKM0edF+DsshAc
tDPCGOf4GPLLw3SjnGMB0H6TIWNbW4PZSOi4nSCdJnNB6bmdo6wzmrg62IKMcerk+n33G0N7YT0/
HO8bmcZLkBs5t99q6iXlkeJyVfAtUcjVMQfmkLHloGD4ghjBOXcNhuWjh2EnWyDIx1j0fZGqHJOX
aE+6oxKf+V0EpCQmAOb7SOaofc+7MML59hkncSty+mOJlLGipJu+nqN1+4wYoHCe4ZMq0aERjb3y
JaeoS12O1bytjG6XiJJnbQX2gcaHj/Fdk+kcoBm7Ah28BaBWB5JR21ABJI+O3XllPaTdBuGj1jcF
7pOWp8gQizuyWvb7TCAxC9lORIC78cJag49BxBCCiDHJtRREv2ZOGLyJupXJwuD9imErNL0UX8f2
Iym6hMojLVTRUQYZLWv/VeZuW0Rz4ik/3aoz9ltl1S0K/zZ9qkJL7kvbv5j+2wNGkbOdLuU7TPDE
ME9L9y59ySBaX8ESblJmHjtogwFp7YGREOPwuGnaUWvA8HuShupw1OwBQgD0hGwmt26RA3PWaFfi
z5d6rmcGrcNN50WwmsYPzKEq6O2mZj59P4BDnCHVEmRiwFYx/GdCtshBPmEu5NzSQ6dVmXyJPq6j
L37UO3ZQsd1CdatGYErLKYZKd6jtq4ie4jG9Nk6KpBhAwpPgQvMyNbxxp/iuYLUcviS4ObI/OeLz
xS60ObfhsxXtHhW7caIM5FNnOeHBuIr0SqhPyT3IrHDRbOUrcdrNaRoAiGiVCzXR5VPHQU6UN5w3
0ubQyyrk3oV450eVGiyBnwwQNpzts//rLCsSXSIz6h6dDXkbny37J8MeWnzcgl4BQx6RQobUi3M5
23hvl5V5eNmVbS/d/34ur6iP8c+FC+GAy6SyDBNy8XfiDSFExXBSSJIKNqoQ0j3E4XbxNgIEeRGn
47jRjvWxWGkzHFte8ZxH6y7ceEYepVPapO/Nbi8iDFb2Zs5XI71RfNsWC/okIN642ojn81lObzpq
WGxyWqK8fDXcxLKzKzLfPxjodv9HE/vCbRI0X/Q+zIMq4JneroxQLyFScgG18ib+N5WbIA9MtbuX
U9sobKt0AqR62sU7VlOfDO2JXDJXkZNo9XrI/cqfb4ZfIuDagt2UBFA1x8TjWhVwbolaT2aU0R46
SmBkdew4OIYmv+B+xaIx28lurwaf+ZuAozDyw2PYsZt+xdMmhrLZ9JwaWiMBpLVwigr99G92TKWl
zUivHZY0OvB0BbVotOPF3R1FRNAG2i4hRjgTZTG/EHsfQ8U+FfcTiQtAzqt9VfNUqMERQ+0B536Z
s/psl3/oJYMYh25KE7Pd2xSxwcFbiKtldO9+aW63SiWFcogjK8oJak8GgQIeA7v41VjonQZSy/Rw
KcdPyslQrzb7gJFwnfVck+1u4OsRAIadAo1KWT278fjKybzZ84N7CSg3WOtytH7t4FxsAKwVT9tZ
ffzwDKQrmgdSnA/XqRQNO6a1g2y+Ys2ayg49jgv4bT/Xc2/ygo6EPqRtt/CUOMsfkq1D/mIVgGfw
Jk1yntpORTbjxq8YJk8+ZYiodeKbT9qQkHOHzBLq38tNYMtXhEGnVFMHpvz3hq+zneEPFZjebsmQ
rmF3t0ryoixvtI8QxCKn/2hDMaNYngOF/bgZ17trRyoBk8C/Aw/XTSF7mn2UmwEUPHjC0m3w9OAe
nnCjSEdspHNDGwVhH3IEzJL0Pst9N+K1JJYzZ/hCrNsNW0+FLwpCE5Ruy2DAVHwfyqipnbdJBYgr
WvTz9hxkT4ObaipMptHXShtft0wqgKgXs0nTZgtn1xc6qH10bmbqA0Ys9x9QjMtkKoR6vzXkweJm
rQ1bvoxz2cZDvw7mGRVSFjfPHFiOvgP2z2OdHpaG1SxS9Jup0seJeZhyVPWoWwPBbhEVIepFnnaa
bwrcrvlK6WfkB641i47jJ7Q1+xruVCiv/nh0COfnszd7REH8Hhm8LN0fpJyFa6GCwGqEWHVixlDf
afNvgPCA4T/PTJqOhlFuCWWzJnCPJNqB+tlpexIqVkCWRa2XcvLakMfxOVnLwMjPGZcw+URK1rGA
1CvCIcZT9b5OzaUqUNpprlXf9xYf/U4c1kL8bKREGO2Zo6MzKk53KGLsBsF5Ovn6XeEhqJOoTf9I
jJOqqFtZAFWK72XYe53DvCcW+cTlzGpGtGqlRqHfhWmHmr6k2QRtY9f/+uWJEJLjkO6pKd8OA98v
4BWXTROQ0WCct1xcg48hOXYe7Uan/lXCnlwHCo3SYC2yedG7uYi+R3zyYLkmrXRuOH1uGhrMPDkF
rDsrkftdJUsaMJTuDV5KCktsx5BsqxJHkqOb3ToNwZyIO5Ek9xNRH5Q3ctO60wvlOBwQbLJAS5iS
OH/fu1+ooBI+Yy0RbX3q99DfrCibYlmD0IojSekZz6c4Ed9J4LUu6Z+HTfk/N+oGydtNdWhwTq4c
3yBdhE0iPV31XQPIQnbNFaynz3GHLAOKmxGkmLKyiwd9kc5Z0NaKkbh9kdkbARguxMh95+tBpZqk
oyM6VvIbpxb3Su3+D9sQJA5R0PvMeSmM3S4F5nUF+A4Vwgm317CCe8Zhfq32HMFiQIFAgwxySSop
I3ZxTkvEdb/6P2i5tCcsszyG8ATHRH69BtVb9pVRpGLESi+q9fSUVM7+us8EN3SVp/Pei10K7PdJ
sPnV6rCfELzgGu5iqWE+gqKG933HXLRybh5cdwf3Ssb4LQ2PbFF6EfWHXZVZKBkbrLRaG+JxyxtE
C3ChUd2Lfb/Sm9z+ieT1JrMgLNr1P7iENjO1f8N8ZuB1OIpXNmp3OcxUwCrcNCI3ZDiZzmuWtOdA
LDR4Wvo/6Oz1JjMgtCaTwhtKqn+oauYuEckhtBSKJt2er7fKpjpOOIfulk91W/03Z7Wj23ZBVBoi
EbWP9Dqg5+aiWhbJ31eRpIFhZnlYU6w+dEYFb7u3eH3MeS1SXDBioW9Fy0n3ZZMnKpVAQCBXXoKv
DQwtdqots5yAaadlG25sphLeUmOOLUs/yPy1lyU0Ji0Bjrq9dr2aprWNMbp2jDxnq7LW3qXoSBdg
S5ioHAjY2myJllJYpgUYhRffhjQQfVviwFdTPoF6cw2OtQgLqguoCxR8lp3A0MsS9YUG/9Gy/NWl
lJ2MmtkLf++DOmZ/tmIX0QuTpLo+c6tG2Y8JFaRCqAhYCfxwVyk4jBMRKlPCSIMmtAX7ib6XiMED
HCOg/L0qhfrEPBMlLzV8Mr3KH4a73EN5xeLNfVIkL9P6hzGkGlsHXmaUA6yGRTTVnGz4Mq9VD60C
gnobi7uQsqdOGKxuRj0JH4NsURJRQeertBJqBQy21aE2jMchNEFWQCUIIGP0DHp9Bt4BbQoQ81Bz
uiL8pKv+HBknaWNb/hZWA3sWa9vGdogKgQjk2MP6yLFN4T6FDUcrhxsPjGBehv/gOP9aMdFcBjtY
M7bu9t/H3wSNlm8Z9MACCzrL98G5+/0Jmp5f3ZKd/g+M8wHmCP6isO+duI4PeEew+ns3f1Roo3d4
fP/FlsYGtB8ILP2K835CPboWeq+05K49B/G0Vn3cjwUItWYj3slCK47ZU8ohg3JEcyHyTstGcI0x
E308fbcQMsX/8tDwl0zpat+E/NpYUbzyLMFp6faetdiV7U/lThiCRdg957EHOxqDrdvO628B2+E3
AOLKhLA/0R4iEAx+323YfJ6VtrNjkHHyXgciwdifZ8Nur4eDVo5MAvfLjO8Wub/QOKiTsWJcrTfH
j4HFEHIrYxWaMqlEliyrIHuIC/wCHZaJffNwuEMHKavFifUA4MCg/ljRZkL11X8NsniQGCjf33AN
MnS9yWtCTZED/Jf5RHl0Np+XK82pb2obQtNg28pW252piYNeaU3fycUb+qK5iaQOEv3KwD4lmZjT
q/pvrkbwGD2lFbXhmqksGheUwZhHrmmhu/YNpLaWMTlI8sdYnWEeB16z8BGLGXXpSokyYTxxlLl+
G2F4Oai9w1PZYCmAgDefPGxmoeJDUerbgnucGoPiiMOjDHNuHQuBgzUmQA5B9z2RVMhCz0MPx//C
tu+gOSLF2zVwuWo+qoBXCfz8zhj0WH6lM4i5ZuIFvAdO2RTeGkxwoVq/sRfoHG3kOhaRNeNbG69m
SR/IKE93pQQY/OOiNKBw2Alx6dqfFnFiD3C98nhuMZp7WhK8YGr7n15/8lUFm2a2SWtH6RkBELwU
IomyO7bQRBduyJhcOrQ1k8zMp4C85vsBsSP+a3GMn3+ZRxvlVQcV2mFmFu0j4XwD5KfPD1OxjDdj
4PFXl1zDE1cPcqWgbTf0ak0IWIQU0KOUvPz/JRmrMbl9hAfJ+uFSvaA8f2jNCMXJm24txwcWRRYs
4MlOHMx5Q/AY8TOZ5ibqfhVu6dFuS6+CCOeg0MLfetMdPn/X0gQt8VFoC8TLgbRA4AwA5EEQTc8a
e1ENynUWNGMvcTRUGMDG2ZLAIT9D4ZCxVF2DzbFH0TAYk3WRO0je1FaHYckluADFt9zPk7eCPsi+
Bt5M+M9oCmgV16tZEHFVuXc0+M7bUnhu5/NWudAGjJkV/FLnNCkPR7FwKjbOCTRm7TBUL2Elgz3O
ZAbcms7Mxf/adHCOvR87Xrq/5JodNiTh2CFmcOTssRd4B3oKLoywbCocSHw3iyF3nZ0fFcSLSDkP
0saru4V2AncSvKkVADf0bYrtTxtZjv0zPM2SE6JDg1BserLnVRMV9pIC/axq5V/oY02X12Lw+zoz
8Q4OA3uEvnKg9/0B5LzrJFWWvEUW9qRiqRoC7C8hVo3DIqnzJMBOjr1SeX6yjY6bqRuf2EKeE5d0
aBCzmd56X+D8u8dW7PfoDeWBUxz1ujsJTaXSpriy5LN5SRHwQy/wk6J0bbBsAiLd8UgN8QY+MpMt
qVv1tfgKh6RfFdWDFSce7ncSnEOFVsdovdNLANMKuQsTFiol1Reut+pQxLrGbQNSpNeF8+fpy43P
fs3JLhQ7GVYjVrK0G8q4LooT8RspfEA/rR6IEQ6PINAKgyKJj0H1t5enYHOuRO2c9njngw3AHNxW
Xrs6lOeo72/HEzlrjYOs5sdxVdLkfS8CaSGhkeVKVwgN0BQRI57GeRvNjJ5TBxMlfDpKnKXAAcGf
4oNP/kYRUxKr/ZCJnD34/HGhDzKhyQeDStjqCfNHgX3Mzudw+HO9WHAJFYRvd5jyFVgJImXSxolg
2nnEg/UNWFH9t8pDmExk96y/zhNlIz9T74rU5pIRZonFetfb4p6rNrmU2s3By+bqF5fj/ELJuQCM
sAdY34HMD7PAwOxxVRxpRLO61F61+2Cs79PRHzucN/Vd6gThF11SaM6Hnzl4smET1atiudIUETgT
ZK8P36jffl1K+DopvA8jpsGnEo1OpaPLTMueHPQrrq2V9sXzMk58135S3qF74QQGyo2fhe6LMWPa
eXU/o3Dyxe3CT+Dt32mnpYV+R8GzKtuwHy+/XjSSJUw0jIiwtNDDf5dMB8yaJFp85vWx3+K9dONd
dBaNKSXVBL2PUJQBHAej3+nwtdyrlnHY0F46MEKh/u/EMuGrsWahfxDsCpU0fRFI935U2z8F5tFs
voWFC6lCiioBMP0VSfyZ2mmzhL850HL3awKhogZJCD4Nur+zehWdT32h6ftA/lL8bmQ8SKI4Lvku
1N8KS2ywidNYL5JoFoDZHtG+CsJPV2rIOjRv2wMrhXpWMg+mIMstWJiwyFxBxuhruHPsfOwZmdPF
grwHqAmRig74TYU9MKHL9wNFpzopaSi1eqkFlGl6HVKrEsZO6eIbLzuJPT4FSIppzNgZAjv3MkS7
UP5uebJa3mZss8bzDcuqn6IWwaLnDf9xVoQ69Ifjr8+Ey0CC4UFt/RS19Uo6dBD/g8fER7wqSiXS
uUDQCwGiA5MCbg2AkmCRh6CxtQgOaCqGVG82hyGS0Izw5V+yOvuwjtSli2P6Lf8/6NydPUz6DG6H
hXk7Xx2o2eGENMeD5Gm1nXvCqnSQqbKtGACqckw9X2Ae0UppugIjKTpN029foDZH11lBTf/M693g
OKTkrk2N3lpCTg4r1J373MBKrpQASeF9fVrLaQ42I6I8WL8UEyzhE/K93NTPhpCfFg315RYcSvcA
t0QNY5kL0ie5xA+9zSnPw3BgfUX/eYfAtpxAREEVxcBwA+Yokry41crFNqnDcHjo/Hvsvd7MIjdk
I2MxpgyxfvmnxYmysUfoJmDgCB47YjKjrh+zsxTyZ5ygizmAa2NvoMIAq4jezeoCwwJLRVZXppPw
o/YOe3N1lqxAHwRLs9TQq3OrJAlxFyq/fXsfotfUL+GuYJ7QA23K68vg7jdWsJDDfAxW8k4d7Sd3
gNC4z47AyVVdINhQQ36qHPc4X1lKZ3cD0fYOFm/wAGfLUW2CaBoa+qi9KG3mfvtE6V4mfPBD4aut
U5thz8kjeanE3NULJmF2/yZQBmhGx/HuZUXWL3IdgkgXuCdMjZkex7z90uyxSa56ghDQt7Q7V1el
2rVp/s2SRHNSq1SXEdyiOpNX/wU6dMaWzBhvtkcnrEQtyPKonB0id4X8BmQIWK+3m0Qyiw6NVZro
ionM2P5y89I5LzC7eUax/g0efOKMB+8sGUhY+1mPjKOf6H/EOzzhzjpQdrADHdYXIRxTyZAOB1zY
TieCPVz07ljZmy7fBzG9k8z8a/KBo1pL1UIGU8+Y1ldG9zkTdhlMVTkQrCG2RXzw6ZXOSLS9Vdmy
eZ3BXOiQ4iTKwqHGa9GrU2G5KJgJYUlAiMw0p22sP0S16aExTH/KNmta7uMMq1qcMe7fMZ2gPkD6
uoT72KoyzeYeKjYfEQPp6hj2511pywaPCkB6sVNvxUbPnaFfrKs888N3rdCt+vKpRiTQk1Eth+af
UenMi6YfqNtsCYac9PelCWir2tT8iWfR9FFZLaJ+x8MpphvNB73th7XJAARuxYplGDaeYBn1nS6q
nnTgra8v2kRbEB221cvvSShnkKWoCDpXceEQWykxTDdyLcA8oQEVEOPtBDztc09ryaTfvY+yt4OF
p5cTziYb7Q7sA7uZJir8RvfnRLCDwwQWPMRQ/hKQI9dCGxefCeRORWJUIJC3AGprabqa5fS9pUEJ
tZr3lxx7ug3dUhwdRO95VOFhbgeCy6/eI7Uk5FxuqqpTjOdvHa3JgzxZFUH0FyqGrw/fWrC0dtMw
4k5OhoG/Wd4iRc0rQWV5XK+2OOxy3sOd7xooXE4eioiH+zGehqIKCfPIwJ1ZZ9E1S0TLOg0psoLE
H2zptuck1AgRQU5xuqFt7iZ1Bfs5AHeKJ/gUSoNMfeAJTQrmUfk4S7cKt5QPN307TZAl6ikHaA4/
xYSZ0UbhN9VrbQ6fWKnmj9cxXE1RXCqgJKga0bo18tLuSpP+cdMWVhmK/KJG5L24Kxx9kZz5yr1a
6HORKHDIDLpAs4mUIsVtWuyQuNxDvSOIhZHqqbJoh/nnURJNPgsa4WKcPliSO2rUl3broKEjP8uC
hetcmM+GkIzhy3rJmWE2XBVe07tJcgfGf7G9NSZx+Kd03aQR/s3wWe9x5UwK3iEMrfPqwJdu0R9X
jTJd3MTMbiyG5FO1ISWTOsLR9pQ5Xhtq7nn6kxbX8GQQEFfBbofxwtP9mbo41Rih5tV73ei+VFAc
DODgrimAOvoYToKNKlHMxgAot0uiqByPAsQ/hxXKSq0xDfEFPac4Yq9n48HY8H5Ba9v+RsXJj1oB
rs5FAOzBy0Mh4Qh76aV1vOocBNdQDpSwmLbei1o5gIVfJKq0Nk1s0XZqO/NZJ1P8GdbwUyxM4bCu
c7+F9EyjX21MvLfGSR0aAZ9MnVHZyyvx1deA5MKNsXNmk3TOECOZ/s12zB7n7XEq/rM0kwpy0Sww
cev3aNW9JdOzOnIPkDOvUey5GOfmtSfsg3wbkcWac3dyOh6tZIiJb7FfOl4rBOWw2HqtshbyDnS4
9I15tS2AQjm5D30f+7kok2h8X4Ypggd75Ejb1cLdmQBBiqSDSy/kXaEI0MbpP7iyczpDcwo8Nz5C
T9qicgvYZEPQH3qLpgll2YoBMVWTj0ctQvg7huYp/3Juu0v/VKaTl33hnSs8C/j6rITqiCitGX6i
uU8CeOZHgnvHBGjsM0/z/V203TalOBravA+9whNxPkDHxvtHVLOq5oAuXQvWvD3gQDocvGnwSZcf
91saFKLAchXwdwE5eY1Tk89AZcAtOD/QFm5cxTLKMEBslJPYtm0Eza0eWROOPIzb3kBQcSDONO0H
sQREGoGtjanT55kBCW1WEzqI54XczA4Am+O0x4pUdVRMmOi9KFoEx2NGg3/Rb+UDl4yqfVQreA5r
lw+BOr8UdddeuhRIfS1ZE8RZN3JC/B9qYahAuxul217oEw7uF3KzZ9ZvYVVqjz/gSDgm9/z5F6Ug
aJZm1BKWfNj5ws2l6xHCTTf1Q0bWm4h3a+2xWbUidip5fdSfxans/ikYBm1sp0hqnQMPLRqK5NHU
HWF0E+yLOOyBAA10MziHFQXKqf5G4Hw03x0r2cF0XryHOx3Whq876cG3li6A6bmXgGfP8j03Sy7P
bGMnbiZ5wNNbj+7XUTjowpmBgJn2kOgW4s6/HQizegbDfo1mqrpiRZyJoijylm4mMTrmit5+pojG
rGu05PJRaGcWoJfJwYVbFUZq7eYbDCvtzHsGrhDAj4KC3Uhw+MNrFiqRzKiveUwS9zeQ2/2p4kfT
6SIwB9Y/mVhsQ4PYLKBAqgFsLN1Rtg73+rRer/ObLWSw/FYnh7fdyliFImpN+FwFKgRGYuShahv4
B9dpBnGwN7JoR7xSq89cInRV/fqdPv/iuhrXbN3kDJeDBaJPJLliFHqxjA3gLM2UYwYGVb/UFlaL
a220PfJ2xvG93c7xv3B6CkuFCeQ1NgUg+pMo22+W404jCIjWkib4HAOctd0syEmCNsNZjgnEGXcf
zmWAQmE1qiiUOxI5OsfRYJeMlY1eMbqh88pFXAYIM8EE/3HiHaalM5vnjlkCRaBpt8a6HBkkIf3Z
0H6wZbWIshUHTG4aLXdEff75zaDNQDz7524CWxLVBOVgqckJEQoRgv+qRsQzhBAu4F2mcV54qOIp
hBdSgeK8BUckp8r0HNlgfY51STo9VyGEo8idzGP5o/phn9L/J2lqxOhhkG5JC1sl5POLhAISGWuc
Ajn1+uLXc2wbrf+0kCRm2+jIpa3U0vyZU1swRv232LMiVyMi42BW1DotEgMiVb0G7+tExKMGME71
tEmknW3ZbybMTYYhcc/zJ+doeyuU1O/J8BF7Yp08qk+GvK+SoU8rFc9Ub8WW9ky+6+ykRxBxFFaC
3sPBfqhprbGYYmgXlZiZsJRXvByRF+9jOBSc7GxY5JLBMuEoQpex2qwJFG3E0Fqp2OCyTWPpdjoX
3WoZH01BwCdPhFgI/5HgQdTrL5EX9nB8pLx21WZUz00jcUHOLoIl+p7Obh+q+UNRqIR1BX9ttEqo
jKj1Ve49w1/YqJKw1OR/E5urFkGZkNfG6E8Ecpr4FCKGNnIPnVuwlQaX7VvBu36WWbJvIWAdt/JE
U+vYAcR+lIsDcMofB4+G4nElGvcQio0j1TQWS9yIY8XBTX2KWquaawuSqPbf3xPOaFuqp3sa0yJe
Usvs1CMtyLfJLpU6ii4JeqYFtLdlYx/kOVM/6R5sAoBSolPBuVzbJ/sspSSjomrbGAbCYPHJoXuL
fXrvwkp6BuEAWIuu5ioEzSbVIfiqh1fVaGsHPqcb/pCVjR+icjDNqp022pZ/7POycTCyIlKBK1Vn
k1yAnHcouQP/2v2ozIxXWG8fR3TalPDN45JgD3EEUAC8wfTRkDZflebL0MTYWM4mTP3F9uq1qM1Q
tqO067l48Uyw/n6eXS1G9LwM/KvYCpBJ4qFuIizvkBGEAiX2mVYZaoA9/WwJiDbdRvGpbjEPhUXv
Z/iF45zZ9fGs4cVBnJyMvqqmXXl2kkgcAlOUnYLPjBGI+H4aTHoCD9XjU//mva/r6jUI3aC56bH0
xEROGk0TdaMcouGTjMoVyP+iS+nNmEf6ptVrq8rEE9+wZx6uDuTnJ6UsJ+gr9C7m7SJnyA/j4eKb
SkfX2ORGFGh1NO0sI89IvR4B535ueNKkgaExaPMZmDcGkqKhpGktjVlwmsAuqI3DtEJx9VOQNGxP
HIo/DjTF5cHOpiXL+MqOlyu2fubBtxMHsUwR01ql+PHTbTv8vjkcgVlOxb3K9wsOjVeAIHVe2oG0
6d9mSRMXERKVD8soiNVMFv3PpsE/ZG8NueLs81G+b3XDHAW/dTMATQUMKkV/dhdqdeChp+1APJ0q
dY9FyaaRjX+Pj5gp3q6RUPnymLrzOybPeIlXQ47KL/LPGFk8W4FFX+CRDc5fmXwf247QtBb0xR0t
SUlDy6eJIvp2lKG6NXQmKNSjzM3UWWb7v6HAvHDPOZroPTjNLwm5QjOWV+c1kGngBNjqNAfciEun
ogqYidgn1/vEzFyR5wuAEEZf6zzYz/XvCwCh/OlYv8gnQnlmf1ra/YDU6E7Op0qwvbRvzbGo39P7
M2B9QNbAv4aqm1U4iYj2HdbQD7jk3NsIxFkGqcTG5QTakA618EjepBXjCN1EVnNvu5phPD+ilMXY
a+bawgx0GwhXurVDHbu2QUQz1WpG1cRnrSIGSdgr0SMtjUpeieiXTargglMj/xoE9N3CEwovEgUF
obj+DyNbWVHjgXsaV0V+9N+CrAP3mYKlvYp+OpQclXbBGo/yYtl3R/SAJcHO0UUpXTAMaK0SBrlr
hI3gIhgiRxKp+EWv9eouAwBOtAuS0s6b4WbCiXnNjO+j0S/CRexTeFWCjEsUGULlIJGUY+xPx2g2
8W8/OuMRXYXrTbuRb88EOMpORcDdbJwO59f+234IdJ1K7+mR+n+4YVFM2w+D0Wk2E4RS3MYK4NG/
NrvYGof+5cZB1ji5smsa0vWW8k6zYQBZa40JmomqxZH6Xh1ezjSd80Uhkkt0j8j8oId3jHsDK2P+
KmtDT28e8vNDAluOTy8YlwKXcrcH9RR8sX/KFYpR2d/JSfhMlTWVyX2wZAUBQFzSn8XCE9c2LtAM
S878T9kFVOLugFHpn9OM6FP9vpO2qiQb6kM6AQvfmwc0VhSHmiywGH0x1vkIegLpnTb5KmqnyyNP
6PfEWqtBAZsBz7sALj1xoy6H4O6o/sK5rJ3IMMXc9Bowtt9BNpuDmtNZmYZuHmhvjc3VfH1nAzog
XZurXzvRI4+CAg05t0lU6K9IXhjrh81SA68CwIUgD9ReOMsnPF+oV7LS6TDNURk1A97YDWws3+dq
tOQLTpKfjLZs5uumi4KEOM7HZJ6Ycnyakn+sBR1RYCpvrfhC6Ap5iq814aTxw7hCIcLLMh52WFyF
mY7iPsVLhvQPkmcEt4+0McdBs92czz2MXhxao77mYBA0JZ7QUVAIXp/TldGnivMVTwwzhe+avhPu
bHexBRY4Gftp+1zm0mJqQaoAoOHOJHpcCr1lJPTzpGTQMHf415nBnSYZCfhh9PbSDJkEalfaOA08
qBv7ysPHxMQ4cCAuTHSXmfP6kdNJNeitaI19C5yiZ7PXg6tVZOXifi9Pf9h/HXeqWFeGXlroqe8E
gUMgvR1WyGiAFY+dtRyS8OkpHKf9QSoXZKhkba/9e07KI9zltwzrvrFyH98s8lBu/VhjfneiPvs9
T0OmkTiGPc/jue6CYF6O9E7I5i2Y1SHrg0IADEg/yuXwsABreKtUyPYrNDj8C/jIQKInN9I2IbDC
fskAEu/QM8raueuvsGE1so/0JTEyrpJJXPSAFCOMLbkP2Fb4HsiAkJW9vbLAoT+1bW98Mc4FnUb0
+2Vxkinh2TDYUO9I/7JWKReyV5PDZ/o8i9h62BTCmNRgW7kOW4Xmrfz7c11pnLfQF1ZuT6ti/ZHA
4D+rBodimpmfAEp6iA2RbxNGQkH2vovj5b17ymaKxq+BRk9Gcire1FY/aT1/6dUzDOna0jFO0Cit
8bD+2W2BMXF8H4Hf7/SRTQ0Or9J2GJUKN85Td5KMgqzjIPnskjKpMnqVn8IyYY0rd42mxIIVA9+E
nCSo9kvoRQY+mMWzyfQCUdGQ5DhdTC+3PBFjsL5IqcIl2M/rFib+yKYyxf03WvHoN6hGlXdiQNDA
8gvACkgHrftJITSFju0sXI668B4vwOJQxweGvsTazJ7b2kAeRWk/ctCfmYkcXix7VNpkYKPnTUlD
vje8uvfHgHpjQXf8KlhhFJp1BtJX15mdzbyP3Pxqk2YNB6l9Ypr+Te5h3wdjZ1EJdqVCrT63FZCl
uSCBaICv4lMxwkJdm+cY/ei21tM+qQB5aBXJrTTymE9ki7Fq/gVGY9uzpKb9H+3YnYekwCUmXyyy
OmHj/n/tAq513dg7HTT+8lwByYS1wHUhwP7s99NnWhujBOegsqwEW0aF6aqMQeR9DTOiR/ZM71l2
Ir4iBbvucZK4Alub7Pc6BnQFROS5udr0XFibQvjVScHzhd/ko9repsOY6+MiVrgoFC3UF+hCg66u
Upu0brd8uPAHb9sy5OAETdHozCCtTF/dcPeEoVG5mlKXAWGfzkNQ6rfyjtRfekPVp5+Ofm60FUHV
n1PjuyH3qksjgLHnpS2+tXEQNrvUTb+SxAe6kN8yXZaek4nuyGxiyVHnlFt2FVgklBaCcTDW2c+x
+jO++LIi9cUACnmB27Mv4Fnvu033PQu4x1/ZgRWkCYJF2ItKxoVNaZQtfV7GBJDXt56DTt9n5bgO
rcCt2EhGbUaDuAOsqLw6E+ptBWzszjpUZENNXJA4QeBR0MZkwnPbI/3RP75OHXVhW9iPX6lOGOQ6
H2S8m2IYkVBtLdAFDqVdhpijgcp0QE37QvF9fUWvGjMnby2tq6grWsETi7CkS57WbH5fFadhDclG
iaUKClStTQuzXtpgn6gr3/z4nUxvALUnBRx/Gzy2m6MxvyHd+sttX2Sy4HHpZA7s0xy2W9gZQ89l
/r9tI8kSsRUQSDKsq2TPeC25V1Yr5AA/iSkuPXDIfgg+HlZnuFoMdy0CkrivGbb8WH+EGDaqyUF0
LJr0WonEChhhvvY1221vYyLonlHlH/R1zDbEiRUxlmjElhC1IidSJZ1590fnTlkY3NTybJetuwWs
1mO7W7d/YnAirMjZwK1iQ4OtlcIfBD//NkiFEAXUBr3QlPJDjReENnsyzkPFjshGeOHqf40VnBkr
KzGqPBm7LSaYeGTXMj5dNC/PeMesQoOaYaFf1TMTjsorlfNMhnQzFJnrUq8Eyy9vw8O8oGrT9EFW
X8GGHKLkCe2xbvhNZgYtIDnye+RET9GMaRzEDSCpm7FBhlkIMaaTrGtr2XTmOXlH60NPh0E76TO5
a7OCXqP2+A6TyOU+mnpN8gbQXxuIvpPcaUXK3Q9VCzYfxgznu4bsjnfVfZewZ8wOeQV7+jbzUt6G
+89/jRE71RSjyZ7GWvUpInkuMublSWUccoa0SLCSg66+uZb8Fc+8tV4/MQOCMlO/nUaoWQsD/x+/
gkyoJiI7gwYjLST88lQTA5hGWx/rDlHjzlLCyEVMHtO3UKB8cjGnV6OEfjr3f1Nr5zEOmK0I0hfS
ZtYVFbZDc4WVAXpFwGtF9PGVfLPrnWeUMcUqMRO+u6Nc1yJGpDu6GvKIwjqjbKEDjTbrSwFTaVSw
SoW9JORsiMhOFYsxDuKNv69mGXG9b5TW/8QDt9btDw7eEqRIpWu7DhBV6zWcj/2jO+NLKJlMkqg7
UP9FZ13yddojkPU2Hfnl/QJ1JTMT6yJFKAyBKZfSojWzh3uAzpendLpXEZ0mxsDIV4f6CKlRCYOF
q9PMb0XhBnyv4kau0zvc7pVogtAZGq3VNA5gxafAvc78LzAmY2tCtJtnK8FljLLa5pBfmNZ/zqNk
NtN2qo8q8DqX9D79+I4aPkIEvyYn2kAhKHDaNFJ6+N1ZB74ccMqoEdLLea2pqUADo9Jq7U32li4V
nqx6GjDlp/H2/IPA0YhEbjoQlxbgaU0R8a6B82rXBpLGF/BKgw6dHT7bu46ReDFYZWJSRJInhhP5
Z7InnYr8PVVvgIKQcvzGTuzHTIiT2US0/BIcOWOkL1aXlXyubyWJfOIceM/8RZyCeQFt8eGcYXAX
MBDzyPWEj+EWGmaOEfb/qatIwr5+A6EVoQzOhDNOVfD6x04XgNa1oOA7Jgy3x2CGx4QYx+Ijc917
RAlBMZgRhOz35l4nxRu2n+FscexyFQ1DM4MC+9fI3+6EfgutpemHqW0aEmDSSN/2MsPdPpMKdWVq
382vSFpuaUsiaCTU6ROcVW7TnLzIOdg7HoQUsJ6Tdjqui7X9S9j1W1UM7SZ3D2EhdKVOXwU+WJkn
lMrn5R5pJR+tIs7AZAffoUCaKZwqsynolDLKq60qFWyw2yxxZnotCTkKVQ8/K+JA8HnqTcsxEoEg
nifNjPV4r2Ojwii2+qOtU1MHjD38qpETU7ke4aXzQ4U90XXQeEyBJP8N2e7BqDSQ6QaMo3iulJIs
81+hV/8AodsJ0nSPdQaFyqllIGPCOxvaCT4sADpQO5KE1wZ6m1um4KVLbWdpkeLiS8E3f44yBKan
dUbde+XTPqFN35gHsaO9+w1Z1UUAOMahFwFuqo/2LxVYAQwDcV7Bk0HJ96uvwqSHJe4izL3pCNMw
ChPHcE1Gj5AM4dPPOTIWbz210glV2xBgyesOx0/nvzd0c7fmsaKpONeb1tpRx5ZxTIzOcqpsyRhc
6v+hMtBnYvnCBiarAt8rcHWH34d2xuONwLtXFkUhNwnXTKhpnC6pHQgKmDwMty6Rcy39pcYmlbIn
O3hEa4DFf4uVvrfrDSTefv92dSnpyb+R+K7Qa3HXUO66cMDUKIWeNMttE5G5uHeTexA4XGxy9iMh
9H2p782UwcLJp4I29aRB1PJpfUOBHiXzRulzLafED6Ndt/dYOmn6g7YcULK4/LQwfi5PyIdZYkgI
VMLxpiM0y5bZFwrhP6pHvVSUBYjiiQ50cgTp7i1j+KF1hyrkWkP1n/Yb2G3fTEn+OCFPuvtawlpZ
Yi7PodEuPWTHcDmi1TaGTJ6m3A7qv5rs7lQu2ZJABUEcOKh6y2cjFjW5Nu2yMwLKUJipJCaDTcHa
fhQ47Qda1KyCMGHirqMEM0mrzmcxBN03Zlkt2+peDkHygTeJvO+PUCPvDWoQCb8u5KUDyDRL3VXL
w0/wvJLmvRdOkIKnvdm01ftKtFhiAsjKZ0QI36EbCrWfIPM0y3no7npGoAfc5dw6zSFbND+ZKu7n
HVXxApnASHN/nscKI1mRFMCsfEWutsIz3Ob7sxbY7bNuL4n3M1ymMuYJykVVhgvNG6vejkRfBM6y
mK1k0ojZQ9AQ/4VASjwyIIOxJ6A9dtQBNmae2QMqJGx51oorzq4cfx1w5EfWVSj9GusGBRG9fAvZ
lxM5OnPc1xHT1ENqxiRHg3MoqXHVBqa9ATkSJwp+P3tneefm0yUXz9sVak0nHhGOrcG2xT/xCtlb
KYn7JZzaoPUGnh+w8lM8QHz1D+smRHx/dBW+7JDxSclGDvuPHujIMiz2Nzw34tGL11vGy2ZHENgV
sWps/Tf9uzxs+LnXAXVN+vttpUelsFlGuM8TUxEYnYodeP1C2oBuPFKJ9lqJtLCJlmZ3trgey+hP
OJo3+ZWt4EuhSitv0E10UvY1xtkso7uaL9L5Kge5Hyu5aCAUX2VF/CLpdhH3RP4tV0ymbDh9bR2x
jhn9L+L5cpeU90dRWIORZOxkp7XvT+6+vUBYomGxAgx3ybj0xtK8vkuJ4yec3MisKwrKuqLsuMQU
boNXHFrYM5AzIrw1W/xTSqZ+kubM0tshXJkM1QTVyDRAOWtHjXFASzhq105DkPyH6WnNW4TfwOUQ
WfUmjNBQ5Rd7BYn2ViFQ/xV2yS/46SEOAPpcM2dPV+oolXNejnu2HaEHsXtqIjoqneWaeVVC9ba8
ilE7uK9MO5zGd2wvST6DQoFoB5a8Py8KZiAaYJX+6ZGGAxhqgPhVtPYodmLUN3iI7xeXcU3PnD53
zlvVcObO6KneVXUK0IL99YKaF/JFu48E14yqpEhiSF+xLAuG/rNRoeHU+hkIYr+8JSoeoYa2fp9n
kNKJF+G0D7vK3c9aILWlbndVnqOOon6rqCmUvi2U9exrg8WbSddIrPiLj+hf67Mb5v6joWSfnJP/
3rstP07/61jE+MdSpe1Hy/boPHfEf45x/FaJaDDAWSU9mgMpYjsUj5x2PsS2Hy8K+kdulajyJdix
BXS6l3BQtm8o4m8Vh+hlFyCicczII6yptIF4TcjX7Q/LA5UmEabmQ7BouWCNlrGsEhjqd8uLl++E
ujKBmIbXXCpTbqXM7iPWwVCsePMToSF9ZVIcxHr1vD9PKlUUlNTwOWbGvSji8a0M+D0KPJlXmvFa
oayonONE44H4PpNwDXWrWr0IX09A9V0R4hndtBfhSYMNt00Sbo4hMx+Hz11c5AuEq16E2uF1sTR3
o4QXaFABJYQllF9KnQSm1J749Tvfj6MduW9tEWabolWJruPEICNHoFCWGwFm5UBXd3Wv4K6UhwTS
QfJ33UvkeF2wjSDj/LdhYMQ38yeVgYbVLCJ6Ze9/NJrVQSWvfo/xPxH/SX0RwTGMh7mqZepaUYVQ
W9pjeAsTnbqeThbRbouvxqWKLpRzaGn6Xxhc9shUZJkFgE6OlEHYj26pdBz17255Mo8yy6TmdWTA
h6RAm3A9sPo/5LqaaIyeFvba01v9w3/zc3VBCPJf3X7nnEBotdDrOI3rks/yH4hkSIKQdKLiksAQ
cygQBH0RCQtih0qj2bwGU/0MF/1/sFKXfrWX80jMfh7xBjaGlyXqbUGEsIMOBRSZqI2MDvjB9Uxn
MBAwIdaCUkPqKMhWyfwry6Dc/iQQohosieIm68+YR9++tGKqiVkooA6AOkdhKr4ojhN/aqk5oNUV
eIsW2Wa2d4UN7iBHGK9LUx4cWuOncTB9X3PFeCtcTYp9en0thU+M7h/8tSk0COwggyAa4QXQ2a7q
2TFVlgXm3sgHydcX+RhikDnhsd8D+it9oBnDnXcW6sgHWA/jUPSasYlLsTh1BYVAAyrPC8lfvpBH
w/+rwBBksRSxSr8g9krfzjXKV7XUEvTa9PPMfrHzobg5vFl4Ml86+GGCbU3EJVCX8cQrUxtueBqf
utli7uxrM46CeR1K6qwGJz+L2s5ThA7ZAAhCy31avUkY6MDPSnx2cVrFBU1ZWLBn1lMFV3WgNzIz
D99y+ybTt/vML9yeD2Ou9PXfY+6x6bKnZVaqADk7DoIHkQdYi2w6hbyh/W7LIg2TCnJRwSCdS23z
aI8ATUBsBM7gJ+BSOI/zMHR7xjkhR0Voah05Q22RzpKBVZDtWCqH+4epM0LQMmiDCsYsG0JZHUiD
/Ui6tGOyW32mVuSR0vwO9al/ZLycJtgWcVH9IjJDpG0t1HVFVsUDhOLB9RPerISrAcEYev/oRuc9
XojmKkQCFCKtBidfr5lrpfSRUcfyo/vrLRnKyaCN0UTSploQvrW4cUZzOR6uahuD5GF0fT5DDu0z
XTPl4Dpr+NDCQJhxPB+jaY9WbCurQ8+RTmzfCj4LzVaH3Wx938omSJcs0JmV0dfuOUAahRAgPKqK
6x7gIbgPerLiCDCNz4xgoAKQKOJhb7M9F4wHoiyVCCnvOFNwkTTvO0zK/YdbaLdire3z3whJR2Z8
BxLULMv4RhK0PmHScOYD+nJLT2HiH8O9ap0wEl2aT1KVksLxEy3C68VavS/NMDjns+4AqoxHAf4c
DrSZd4D5dCYe7bxSPbPxwIDYehjc8uM82LJEj6X6zxQKTylYyew8IhdCgSZFTzRQ+IqAD/kACxny
/jGmE+DNoqdn5iENMKWvKvWI7vmpWSWpv0nzSL8WNxbI8m7c5OszexhC6PtPvbB13njWbk9qDFwJ
6F02wyhQorslI90qWoVWLUHh/aL7doGKCqXHnUbYacmHILPyd4jlzb6EEZCZ6RU7OOpYITqsSeZl
zDsVbWT+IwkHlPlWLvHszvTC9NJDBTvRRKRkAo0zqH1po1RcOlX2Uumysc5+sONlg0vHfw9OruLd
9pCF6NkVZjWwk0W8qCVGBErfeeGVg622EHGsCSd0/twK0NGAzsPX2NZCZ8y+yWTUgchK6M9TDQeV
qNMzgagP+Z2wKcF0KIuUHVX/mcUCTVwWfTbN8flxjgMmJDIrge8l9p1vNpUxCuwuShPytZYzOqiD
DNmpA5rMP+bneccXz13cj4O/kAfaNJknxSn61XF3ldd+LFFMirgcmvzNM7ZmjiriITMgrv6zDy0p
hLa/Iwu4Qsq4FVkrNSn44NC0dGRphn9BH7qEfEFn5wVagGFRPIO46o2D3AG7Qis17NTyWR4SLBfd
On6JOmyqh3dEQSWdP3calSF4Xx2IxhJZuoXbXsHwPxByk/Ym9yazPDeMBPiAEfkDHoP87lXXKhoI
Ibwlbl0AjOQameVJibZ8uoXVs82nKtRoJogsPMil2E9LnaNilCbMWVIwHjWuR9ddXwf1KNITl69O
HojxcDdu8xCcOxGYhwPmbfrkTtQxaRItDCREHJ0ixHWKuHNhp0NzAJQDtD5GI/J75CWxxH0Lxdsz
aV1GvfVB2HxSRfOAGdt1Ez+AxobDpheG7HC1lqPM02J5C36xO4q8Ns0Y1IfhVeuxPM+A12xujCmV
cOfA+tw2dTdw3ow6kD/Fv4aku/uDgbyqJU5C7q3x3vEpWoEXfHJQchECjsPQEnGTVFoBlJc4o4Ww
6XK/+7CymO/cVAj78LoxxEeEDM1ZQD7tp3xwzqSzMw/wGknm/SOn/xQzJ7FXqd80saLogrYzwupD
Ei4DSLGUCjRw+ptLrq6TQFrJKhY4KTCAk5sQjxNtDmJfwGqTS6t3hxqSU+p/zl3zFm5ruDBzlh0x
/n+qlkorGWeeBXbhJfagqf3kW3gwm0L1HUS63bH0w+9FsyPJMQ/2P1U/1GsIkcTQGpwqriVtydUf
wk3Y6IBlyEkLJ91GaC9mOxWgTlMGTcMmTW2NpkiuM2SP0Ks5Xo/VBYHo1f8iGElhi4fsdVhS7WD7
5NHzmJFfaR5zBrNmVp+rS5yGK1FevOEHe65KsJrhUkcatwHeN8EDzamW0MuDc1orNTSUQino4x/v
wbFkiTHLQa22P7qEsYFnMC67tmd+7kE8jbq8uMC6/mLgirNOav22e4fEXfHcNyVNVFrJDkL/YVir
VxG8ylGlEUUuKETTR6vdT0Ba2NIIaOjhPlT0Axrax4B1Al1eW4ukinKEYugecNUbgOLia2IwW4Kb
/b4QccFbHOziSCddTEgB2uzCLJLuP0EYFkwDsyUjwtYdTonDa8M5YX/dMG3EG/LJYO9vvNcK2e4x
MTerH86upkJWBmBYTAZT7oJXL0SohPpnJ7DVb3MWXE72jlOfbRu5RTc61q8ZChjFUYFSg8ifCcIn
ERo0tMgmmxqizf/9Ho+MnJtSNhifsvs5y04vhd4P6bLJFw1ZbfIp+/tJW3R9Qa6LLzltr/A63pkx
/P2VmE+0vj5If3Ww73xhkraVy0RNMtmnPLLZsz5ot0W+GbTe5NF69l/OV5wjdxH4Xku4kBbE+yMl
u+hd1WslLYUF/VEMe9GwycKeZol+chhI4fEH4dGiqBXXZUU2pnWsOppjA/ZrMQPn4RhxtR7g53EV
sT5BPo6VmjNU2kyESDcq+sS1lvTszS8PHDckE2MrjA2BqZjNRpb60TR+IS9LtTA9jZHEM3uKHOPO
JiwrearZxFCmI+6MZl6DBO1SsE+OmTtdRMQksRPT2yiZMRW/wXcn2qtJcg9yKSQWEM4dmQKtw2f/
CZaRvgiMgN9NdkFrfEURiPw2Kpar3T9kRBCs20oYjVlEnAqzfxavnCb6vXHlkX2Iq2FtKgxi9xyS
yhJWzUfKmEl55wmxR+xkJEScVUQAcOw66UmHyKhBdrixAp2y7l3sqv/7ApUoNALXsAuB1x15L95I
BHLzFlAC9fkqRS1xFUcsIk1ubadurMmz4Leq9aHr4T9GZn91Mee/U1n4HCAVJD2JfxGfm1qWOiZa
bVOIM0zBLyXcq0uFX7gEjTeqoYZlo6xP+0Y1w+2KIy8Gdg+WcvTbQiQShj5tG78n9m4LT/5qtdAr
vBJHko9UFMrJkFTTvDOVz1ud7oU3OTiLw/c8LcipUeje9q0IsNrrT6WOueRrJyxziRExPJ2z0J2c
ljin86dD8hu5JCY8u/yNeTOAkZXB3P1mAdwKnVaBrzyXZ+8GG/DgvSXfbovMuVf4Y9MSHcl0V3rA
bH5gOq3HuNP2I1xjBltZDl6umPLDWhdU1u/TmG/JKrb+tNnrQTwTSGfVIcBLekAPjWDF4kw0YNoL
gOzIrIvC+srB7eKDrWJ7lmHDw/0XKmb+GzX7mr2FtORE8qHLGZFkAqaLD3EfNIbfidWLl1ZC8mcd
5iYfbzU2NGOSJ11+YrUs9LZF1B/aLRp80xUFsSBRSE15EbzifjOv9OVBsasi+0XBFL3HQBeI0z2x
ipMEQvnQ5ss3HHg9iJ1AxZDMubdYpg5LmfnFlHsiYBFgjYpUHaB49p015ol5UJBEc+7hoSt6xnJ6
QBcxopAiqy6FMHgE6yjRPoXJirgTAK4jf9Pk7ps+pnAW3TzVAvdIg2S5+FTPhQUO1/Ypgjkq9ehY
4jDVEfWibZZXhZreD2VIYOLAfxE+Q5xjY8CC4tH61+NfJRMwwE9iXW7MVU7enmKy1FC1jYbbUfem
ANYwfuiltUcyG2o743s3WUWcjLZjgNX8ZEyGnpEkIVxWkxCKFXf4wz+oTgUYgS28SR9noQVLe9Cc
MMHt/bXUZOoazDw43lm25fEi8yu0wHRoAT7hgMi0u+kU/aejFbPRzHAfN7rFEfSc3hybW2tXhH1v
YfdzQIUHGlUopCtc+/w1tOhs+IHkyIwqr/8whuD32xw+hu4+OSrgrR0owUMX4W9zDcXTYHQqYjJ1
rvc39Ewk0Nh6FpZpI6AmJuL/2qt72PreDMn/aJKna8lOB+tl7Kg5+gyApsdqOxiuqe9MIL+SED2B
v9Hbz66ysVQKMBRmmxpJRI76EmZtG11SPb8W14xxZxGGMuz3514BatzHCfLqxyniAZPn0YJLnHqp
fJiRN9/vlEqQFvKQcM7cXRh1WbuR5WoPucw3e4IKGY1iFXnIBUlg5QNZ/wSBFBYMbiZ6HAb0b1Vx
sYViMydGPmJH6bMmNIh/Uq+NBITjetsA+6iDshzed/v3u1/f+qkzThBRGhhQrAvG6N8altlxP2Iq
fTeJfD201knIcNHMesjpQhSfuEFhGkSIKxaHobcU1de501DCU0icgAUqXTn27a3LNkYg6bt2We6E
UUJw1c2pxzk/bYgDolUETfVx8kYlJOmyEkSddkOR0GBjVj6yDNWyOybaZQ/yUFFXfrGvr/fV9vtl
UlwMIkAkK4Mj2rsC5iTk9FdF2waP31s/vpT6ZU8dMTwmbPmtC1JkBn0BnP4KupplpWCtV4dIRJmQ
xwWxm2O1CB5kdmyHAtC7VvPXGeIXLUmaZdJp8uDQAQdha9C2kJKkFSH8UodRaBJR79morGDznt3x
KAok4VU/fyTQnJbQCxrtbP6SsEuKAm9h5JD1DPPY6IcxbchxQAzPRvTieHnqPfCtdQ/2Ik4Lbfm/
UJ2KP2ULSbyhUVIjv+phgejE5dmi9cDyMuBcjWl6+Yb40qB0PX0hv/tC4mpe9OSujVYhbd4mjoEj
GIJdvOfTyMMllwpOG3oXyvnXgc8slFdwacUmrKllLLmN4JohfK+4vIwjAVqNlPh5uZJcdevIXBr4
58o1ue3MXbZ/4NvmZtlFWNb0k9OE0sijpq9gmdOGtTTdPc8KLhNqLsLPWvQxjrGmas7cqVfW+4Tp
JN6sjrT3dLV47t2381IIyRl2uDtVU6qQFE1ZJ+mkkJVeh7qWh5ZRP1l8NuUI7YfQ2QHPltXEL7a/
+aFYt60XIt2q2yCEBANjWcVJuUwkwQen9ZLLo826+jHFmmpboS1EdWQwxsQSFzLNBj1ujOtG5x61
yLXWSwN8MjFBPSnJrmfrCG4wPvjEczhtcHdmApstq8s3wk1qwwkVEl0lbmF7FySNBbXRvbKdNOA7
ryxQZdHQCYDdgxXsQKbyRfxhal1vUUKl0Cdg0uJjBoQMW3OZRX3xel75smY13RCzKzlMRt8abYS8
EkMWOJFK0FZqQ7PA971Q3sAJGHiJs3cHxfXzOAuEbfrwdhg+/Ej8wFSbRfRwD4cCCslhX2Ig7Lp0
gItsEshXSbNB4UwLiThPdByiKI2Etav8ikT5XVjRYDpCaD9NpKFCEEINmIe3YVnIBfUDIdCzEPKZ
/1JiWxiRG3qK3x3WL7iRheQP8Im0b/nLRyHEQk4f/XUBcShAFUYSjEQAZpeCHYfuWTx/Rhp4CBlT
UO27g7+uDlyZoVqQmgBh9bY0UjtIttg27PB771uTLojqB33HmY6NzStXmMjwSQKMEgXbKks0DSJM
anN9DzD+p60krAGjZPatuVCmIy2wsn4zB+etcFoAm7KiJP7AvCTkyeQMsdGLcbTmW78QMAbgqsMh
pCghuYEx+/jKoPb9dQUAUbVKkxRtfUC8PC0AYP1Cnp/0c7Q1yoD5wbbd9UyaO2BRXXN+tnmsd3ph
SLXnolOfYlGsn5S6W10KaNRhAJx+5h8aR1htsbWrivjg99smRd1JGv4yQ8yOr0ag7TYy5hq/l2j5
RG9PPmSe/3po+UynLF3yXcUCz5H5hPngEcN+gokcdWe3w/Po9ubH6GNkIhgxZ91QS49DrwxFh5qL
8agmht+MuN5LQCQl7i8sw7UFSAn5mZEHNiU7PO6YtAsui5Uuugur2e3a5CpAryAWuYrlCTXjC5SF
H/OXAVPfFf8zzGG5qysWc4SJxZN/MiADkpR+eiiGlypazf37Skq920DtQoF9XIGUqnMluiVo7rAK
oJg1DHSmHc8nCO+xmFxxqR7UH068+Jro+wwUYDQBdAhW0KHLRlkSmI4hfoM7xtSWf81Zxs7/ZAhu
IJi8xGGE10TJp2ZeKDiS5E/eHB47qlk+GbofEn+mJWWtMiTh6snU05WCXQ/yRJdWrhdHIhzS4ri2
i1K7ibegnu524l4xdVZTWpazqYKvKC7IOgrnAaU6vuaWON/uXGVoF0mt6uJL5CAXlnQjP03k0yZu
kpw+JDdeUT50lcaTYAo4UyRo/ytJAU4ckkxTXrCS+STtHslV81OYuL5bKlbSQUL1EAJXbM2ew/f4
J+bC31vDfCaQ7Q/M1hlUlZ9BsMIv1/g1jSOVqq7m8WtJZvO3CQ5ZC8DJFqT2se7NPI2GhIjfBNV5
r8W97vK+4gT78OOfFkovGG+sRsyFquDoNI5S26TIy2wv3Icm4A+5FPFapPV4UsfqO0vT3irYxsdA
ddSXTlT6F7F6yyjFpMM0U+JVPaqRtdXwy108k6l14RMspPxheTH5V7Y+3liv/BiMC+k5iBAREe34
sHXN5aKE236SfgvRFzfLZR7FH47C/iIuUVz58G2WQWjHAoD6kcTk4XDOLeJOSa3E5eNU8zmfUHZA
u18b81jpv0Tdz6783ZV9RyOOhMLyVRhkBurIenbpEBqPBTGwxH9mU8z6fqlKuctpdh/9VpSzobu4
2mOvRHu7viAJUxU+JxVCbI/UBJRHfGdC6gnYHpBX+G4EZ6mEWwSDfWUixb+aPjIpswfXdzFTtH2A
uNOLmp5dbCo+uMR+dAWzJg8w3tWgtG5xkfRaiA9uHNhP5VLAf2zCgNxvyRAMPsGFC+EOCKptUb8v
iZDK+w6VZ0gMUjvFksBf+v1STT7p7Su3xSX08+vFpcz9CMsTdBKEI17BK2spkn6jVLEu8NNeW4ud
/XD+vdquqB5msubVz+g2ANWEHx911+dPROM2qiziCEowwSXrpDvdoSV5M3pv9FZUM+x3JquPVsRS
CZafRpI6lM7HHA1wSUk6Rj3u7eq4oOVrSopxlxq/2fWERFD8xlL1zZvOnf68fN0aTGT431+NJpKx
QVWAnWwf3NUCW6U1eSXcWr0RKrvixETjgfcwxBLt6vBLfyLqIH+9NnxqRmfrG1toYMSAiHQM4HJY
hPMH06NhAQhUiYc353cEnDb+RyxoJGTPWYSDLUVLwh9sGENYzLy/4ph3hF0iT23GdK1CKoKAbyRu
aACuKH3IDnpW29+Ckz42naV2yxS6BodMHUx7wkpHHz2/i7vcxUhvec0VKOuw4JjJdZLAsOnDSU0O
WGlj2dVMoVeagYAUwJfn7c7+C5aPTleNyQ5BwpJzKAMfuwS+V3BKgGZDFtmurlUws1FUgeDsW9w2
/9wcHJe5KXvx9TSrc8UJJGcTkvdLjLXMCqC2Ek2K5REH/yjv5Y57FZlY9jwsobXGX3axUZ27cv5q
DSlgShu+ReB7qw9HEic5j3az3s19OtznZqdRh/aRDDawW3q6E1FDvW5Gm0vWxEjy+27L1JbjyBxo
YqhWBf96AMQRjF7u0bzuC91t7sJiLV1oLEPJcUT7tjJ2GegU3GXVZxgt3StezlfhZN1TSXdd3esx
BbbL+/vRFrx9DoP/tncEmO+PTOqMcq/PqqGN/v3eY5qtjaUvM9Sxvtlu87MCMxQ+cO2J0FMSm8AB
MNHZFUlV+5SRGixPgB7hpuJYRxSw0urYiAEzP2eOgak1et8etwUqEHm32W9BC9UqMEZ7Gl/zRPAO
ZayST9oKzy0esSm9ba0dlBE271iNQMpirD6IrDni8HOpMKKV4fgRGYIDsPFAjfQGD2r9soXPCIVz
JEDiIW91NKOGHlOOkCP4CqbNO1Wn30MXd0J8bKPe5RHnN+EFXnKLvcXIOjQxUQjYouwy5iyFns9N
hP5BhCETqs8hS9fFn5Xrk2025GEPkcPQjrngj3hJ0eYiOLKVKRVpKx6y3rKYS3U8yPBoiexiJC3y
ul8J0MHZm8swkItK7jlEdIN/9IyKBTmt1oMhp8lm5jkf3lzeIzhb1h48OHGKyEc/nuplOM4knhXv
TwxP3UCOrE8oacskuGYrXTZI8qbWHxqiE4cFFIGV8RwmuGDQPw1JOYUCZnskxuzK3iKZs30AeDSB
suHENiEGazhrjrHgT7gzNuMpQoJXIVb3GwErjZ+xohVJ3Yzg5OJJQGdOlYOcpKqqSuoMjUoShKV2
iwknWDkh4jnLnrF8PpbKYiP0TILU4XZmWX/JNcYux6MjTgzVLm1Zvov8q1Cf8U5qT8UQK/oynUbl
41her32yDHeas7kvN6SH1Z7PwZsFiPXotOZSI/kY3xgrCxksa7+tYzyUsqXHzq72FCwIkndAuy0e
ekdo/7WuFzJir6L5xOuLgomJgyxjwitT2NvEeK2IIjEAs6Ln7flLeZTTKNqYllX2QxxPfHO8rIpD
liCSxNxv0PMAuYKJt6lAleSNh3hNBkDE1+e0xezfgrNHhXrUW42nVmM5kSvVnV8bo5E+5klC2l4f
tkC7TnKnP1n3ctD7wtNhIEn21Nb59n3UuKEUK2ouGiP3FwnCe39vMhjdGUobMBDoEUzyrZ5Ry038
PgFwL1+LwfNlpm+g4xE3bNQyIVh+jgrMevrM1gRC9A5hgQENPDQvM+1FFNutWZ8b5r02c5gCQSzC
ZoGF01j4R4bFOJomAaVrGZvTkn6NAGoGWvtjHtDxZsLZ1P4OvL9S5nF6v5wctXqbVtVH/OkEOoaH
mjJvFxwwa9XWL3IKDh7W2w3nrscPO0QDxi/Ez2/CcWmSO+kCb8o/aZG1+vOBm2Iffjghyt/u0dll
3bCRZZIjLnB4+GrqqCFZYu+CfElvghdBK9/AN6d5YTKX2C9aYPt1LI9uD34yR/3pGtNBYbosQ2xf
wX9mWfJA4IxoAA7NL8Vt5YOc9uceuEj68whmCTowD/0aqN7B0u2JrxSBUqhrKhWtwrzjcz3zRLkX
2WuNg+LtIoLuzMiC0Ng5Bqd4r5WUp6Mi4RrxdKdBl6UNx7iHrqedjSZszgcilQlJ5Pk372TwFoZc
eFEmRBebcT706eyrqf2wyoTzf0EV1OIjUD/AyI/rP3LGXha37YpBxG/paKOtzU5HfHaldbH2fLiu
GQDvosQ4fl0Sxm0IJPNMSd7kj7aZLdvIEH6ikVfGSJQGVf3SEq97fRHJStFTmhRzmOANf/cpYt3c
9nkpGA/KAYo+myk5+vqDN6whCYFmqHdIKD2zOwR4b1En/fCyVwfs1FaYhEolI0FOpRwhEJAWXAz3
wSi7D2yvbEQ/w6JzghWyFb/5AqumK+H/3wQXs2lVpG59PSEY26BqfNR3r8vE1M3Lxh+i4lgMdI8d
Lmg7h5jdY0RnipmhyssLgsiEs3J4+tOG8PUQ79beN4K3+uMoiAz4k+2lNjZuLe+EERERz21RQuY/
Eza2O/iRq/zDqmLf6+8CqgTtsh0nnxSP/I+noPXo0NC2ve2jNx4TqcQlHK3yUzROw25tZurR4VEz
j2GfwqeopnVXHbfI3OFhia+zlrBpqJQWLLLx2+q5r6PT2RXkG9ya4E4Nr8g37RXQge+zafx5Y8G7
kV//p9M879nokgILQDqoXCsL08Whs3w0+Pc9mKecEf+uFhYrGAE+5i81AZE2UKvrxfa7Y1RWeoTQ
61G4EkCjt0dp6ZrrF4HW393PXXfZUjANmyNR27rpsQRCvkqZBKy804UDausecSLxx8ysLK/CI4SN
W4Khts8knsD7C1q0HXh9clQ3lBDGCP8ZGsgbHp0Sr1tqYlIwNepzAWZrprsOWUcDAxL6jwfr2TEK
sct5FHE7N7MtXWL6SfZSwZY+dSRJ7WILslfuzyOzZWoddt+Ylp98STgRWSoxZtmtjfDIfh2AvLcl
WuzXC5i0FCdJTtwmfe92Ixs/6b4iErtyzVrC86wqtWLczEapWXeswt7XwENLvgsFgDODoNttZYYX
duzQl3KKYSzToNiYphMoS0jJ60zQJUEkYRuYulkXAcsLradtm1typGf+X29WdC6DoiIkzkG8hyBT
gpbCliuu/5tmoTe69jd9BajSBAGpnvAwTL8RJuS6l7iPuj+GYbS5gqqzgVqEzD3HQ0Tl9cUIbv7B
9V1DT0OTy3+fxJUsqq+dbEpIcWoMwlD2UtuFCgoMGF7lsz/afv0yInfganREgNupH0+QjgD2czVI
vqhfBJWaCYVwZOV+sxlQF0Htfl0tHSdrvxF4WIiPXtvx3t7lEZGlTKb6DofEzaflXnf5ZDkYbz8L
t/xJQN+LPmhQaDggL4xkZQWXgp+cRfT3J7UnJsvuA9mok31xh3wHsjsWHCHLHOVcfRSNVtEzM1jR
rHgi2OGTO+OUsnHQo0ybU9eBgVhnoJ3b29phcwxke3I5H6ml9tSRX/sHcYHt479avzi7DYyIqzMj
pTgTA5Vi6jSdyWNVH4PyIcNIhO1iYg3BmJcZp4iURDzMbtncvy3YViashENgpyXs4CyXliA4zP/A
92nyml7G5tKvy1TGx6Q/SogCMLwU94z6Hr/GXwg2a0y6PxPggx2EhJlIkW75cVwpb7UqZXLkMDzw
4nS0PPJHJwZThEz1smg4J5BA8OioIMiWsyUsTT8n2zv8qJXSRJ+ZgvcA10Q+EknD6teBthvbr7be
4KHK7LjQ1CwglkdYQcSxhcgUoRbPD/TIZVZo4BxafyGpm/ps1GtJs+iJ9YAthtPPos2H8sFbOp8V
O0Irykj7KpZACqO4eM9H2O5KellvBEDrTNXCVVBUAVOFHD/AG7gFOtTyGzMSXVtBGcXBY/PLFBXh
AZGxQTG8SwvZ7c5+KDlEU5X59wxtl8b1g5TFqoduyjvf8GJojXkMAV4hSv9pnoecINOZwRa+aG/F
rdlPBRY+2jEGLfHwugaAeZgaZcmMyI/ICUSbn9jW5CyK8lOyQVIoA32nrQebCMQSGMm2jfQ6OXCu
8sU95gOFVWw8QzyGMNTiawaIYcvHmjIXPsSw/+6N0gLHlQywc6ElXpsruADKy0C3ZelSt2fZYa5X
JKsb+OFzz6YFcdVsRRyNgA8yxp0VVXObL3cZKDeDRniMJYfLgQ+q+L6CzhuW4CjnaS6JDrHKQOVC
qp1LbLbyMpgiwYE9HIrkqR2GGVgGfHqURDaTjeYW+OMAZhObXJQ4F7rao9RPfhpAqxnnXqGnwtg+
LJb4SAjFACmtzip9D2VJwthN6U5sRqIVOoOXTDoLQ9iq+v+z3Z3yDAXqV9bLDdSf2hRQPX0UTdU9
+p7ntXajq21gA2rOMhJMvtCwyqIS5EUMBXMmgjUFGbvGJbVgGj1YN1s+YspOqqH3LFCxMINK8u+E
THzg8r75Ec+8ULU8ngpQRkDJ0AOY6ezAl57xA3i06n6FFxwobhwMTIEtw3h8n++CkkAMTzRVBmph
40Im3bjgQrGFx4lpPxYo0BMqkGt59xqZ3utfzgL45GRot6VgmJTVazV29QQT5YUQRXJR2JWK42DV
p5rp7FP9XxRXEbU69gm+TEPG6v0NFtiw61a34HX2540ElWkaHKF2kBsyE+YammymhJhAy8OCXNIL
EDayM5I3urKrwusybC+34tOZ4pfUPAlr6fVJ8GZ/MHeZZZv3fmNBMvqEFKXfhTnJAxneYjuA9GnS
nbrjQ4H+/Dd84DePuiOjvg5RRVrO9WTlQXm5GoWVJsbUvbqXA4rnaBW0R/131zue1mQXjvrpeRGA
0KXkGTYyI2ciXbxo2Lz4N0ctBLVixidmio68h1B1wMHp4APRQ8j3rbgIqbzNmqCqHFXDPw28TecB
4pwIhxAG7l3QCMWuYm2YDl7M4w5gU8w5Me4iauynjjcibKTWeJ3KJqZt829nWG4oymeKo6RGS+Zk
ufzVJ7ks21AO8ztd5Pql0hUuwQ6Rb9JMFxo5aOxe+89ZIFpsrfAFXNo7qlEJMDINs4EfXLxpgdpm
cv93howKCyBTkUljQPsoyw8ZaBqglJkQ0zy/ZC45b2R2mo1mIJa1smrUGS8yLPkjGNZYlNJZhE6O
YugUeyHpS3xHQXiXVccBKiKLJ7djS+eS6KYLTsUPKgu+0gHOtfTNIUBL4qZwbvD5pnWPBvVwaugS
NsAWVlgU6DHgEIgLKGcXK0mG6Jczwt/1k+Lmc7pLfDIlTd4uca/ChyTmki81AhnggoGiZnqpeqaN
ffsmntuecBvcXzbWXPlATstcHskJI4lelc+3TvxXS5NStqcID2EuCVwNjZ/tukUAt2kQO6JhatGv
AOCvKAUsj0tgm0vh5W0KUgehn0sX9oC0/3PxccVnmyMQ7f9FlUDlaDItAWcbEeAKFH5w6PeEs81e
mJmPqN2Ufw6fyNFx5CI5ggog84l/bYmh0Kv4A9W3VhQKMKSTQHpBFLH/sJ17rNiyPbe8EXcGYCd8
RsbbUwIr04S5PbNzkF+1XMH6fSsn+k+7QVrZwwdhCpyat+4O7BT91ZgYtIORWDNLbXB45fNGWKE5
9oU3eYZQmvV3JOZ5KPoOyUJhggXD2PNwUHYMCdd+VDcPi1CBm+kgib+I9Obsj8tSi9PuEHVd3nYW
Ysz/0VXlUt2HycxIUXSmo+bOXgNNmvFIX/AP7/fMseUqBk1uCliDk9pIiL+NT2kDwbbbNBzUyLWn
HbIEIfCCJOvcE+KbdQ8DV+9xWUyU5LVcWckP5Ag7tiv+PaclqC8gvRWPc7V7pFCS6vI/xGnFX8w6
ppSNSQTEHWM/09KHnpSLEgpDc6nhOz5xO1kMaLc+VLQLirHjPO7CwVnsmMI1nNUrrWbc+jnKV/iq
LirMtC+DEdBXgPzwkTW47ZSV0clx4ZheMlZ+Z78qHEDG1jyztanTL8IljpeQwu42a2XZnSx8+gnI
yMHR0LtGK5zzBtG+8oMWH2BhMETruBn2jETU2wB+4nBMK/eecO5klLwelZHaom3TJvM/7RTtLTb6
kpD664gS/5XebIYD0Rs1A4NfeQs8YFVfledfnlm+Ie/U8EMrENjbGTcjGk+XIl1reCH8GcXRz0Bu
tdZWsdltHEo5uuZd2OAYXPiYLVQm25i18u5AYbUx+jEyzgPD4MQcE1tkFZOtVPIsX4FHdgWxfzio
hTUT1SPkpEm16LfROsouHYZ3JyaB6RMyIaRB8bXQrxyxdiZf0t7SPQLeEieetgZaGoc/G3ABk1xd
FlKavchaQ9FOnY2QuweeGDf4sEorEdud6bYKGiwT8tyqxMK/Fyw6IauOPSqSlyLM21cinemNT7pS
1z6i+IrxPEaiYB5aZCWKG41ern0L7tlxScWkO7Z58sXCarFN7dCJBoBetLEQaaZR5LNOlnNwBbDY
z9yXnkWgGLon9PABAovSCQEyauJwzzPSD7m0taJHhwn5bgPUbUjxIFHoaBc8SK5qyjPf2dDEzOw9
p5y/czY4xMh2guzyaN3h36t69qwXCEYncppNNC+dIJw01eodzKpFaliCjs7VDH/jEO9hq3UwtAEr
xmmyqNWTILcb7Q7HpWwUYYqM4xu9/zX8iplRekNdg5/Bf4ZTtL5gnjJaskdkDWwcj5Uv9Nj/qsIn
E794oKNAZk6vDKqCHsZSGZLYBN38SjAsoB7Yw3/fVNmJuCpnuGlwU44unyhR/DZ0Zr2iMP50cNp+
bYALkcDktsSA3tpw3IwZQ1faIsNRAcxhPoea9hvxQqxS6UjgtKmAA4Q+BN+M6j1EFcdauVV704fY
YAChSjruFYndqi7FV9uNiELsrdu46bA4gmoBgfAFSxp78+VcYHEIKuGyE7hDtfR6Di0yiuQNHYHI
xCacaCWiNPx/Cu5AHI3o4BZ6faW2LDf8mQFUCeTC55GfXOSb8wR3BsqWew35qAeUPwxkr2yBNI5B
SbE/8hlBNRL4uhVFoh6FI6lFhiux9ZVUqOcknQV6JoXWG95XnIQNX1spiTxfLomIOl7Tw6FuOuQJ
btbtOwCDAO1TSgPq9bRWvEj9M6XdbaKNRfqp9MLNg5X3IwktvxQXAoAaFRD0FKFbeAnoVlW3ne1Y
7d6RfFMaRBb7hO4SJQDYTf09js3gtadn04kAV/fLRfvWsl0x0vf9E1LdNyRQMN1YtoTf4WkoDBeU
Frez/9rKIkiCplNM79KQNPibb4zXhRJZqFCo9Qf69/qwN9Mxgbsm7IxBTjlRGcmIidinLFTJn1e6
3YNjPsCmY+NbNt5yWgbkYVOsxUyXvXdoEaclUrjpROePGZCoZOCejKlv+kYdMPciWgmxDaSfovo1
FyLAMDBP7ciDVpwOiLnsOgWRW/n4S6Iv9a6E8bq+zLqQmDMUo7s3pN//1gtMwkWEMM3Zgs95s9JA
eRmSJH4Us1fVGquRYrsYHfpe+wIMRwpdBkmcomYoP3Se7lAWHapomAhoYieO0xs1mMVN8FJMUDWG
KR6C+asoU60FCa6BmAx3eoAXFuW+AsJ9XamR5M/TYstoAtjAStJzE1ASIPxo6wGhJpfn7iy3vguU
QFk/s/jx+CgGAybgSjwojbBS5S6K6lyTzeuE7QEU32++nGk/CFcLlFrr1esozbneW64ySsGz/e62
6C2YZzgmhsJazCNkYdRgjzsdQYdfBUikZdB9c4tXpkMqjdxy+kBFMEuvk+Cx55foGQVXxEVJV9mq
zOwqlB0W9sBJOU5p7xhsibw5JS5wjGD1arRIUdRRg7sPhYEj1kcpbLFY9QRRywS7cpKdx0HAn8Br
8mVKYOrO4QFfwikg+6NDoh+7Tc+YBPTu+jesMAbVdVmrQBmIXQvEYobrGjDe2Kca26a+wDhuAbi0
nwkD6508YUbCpxr89JX0t6FAIO9bsMKE8wqSaVatf4FaJtvKg3p6dbYeX1uuulpD/YQFKVr2QfTs
6ubtXA+/rmXV/50q4YbBJfdRyOOfbCvVcMkLPsIwLWxD9lnWL/QJrAlTWz6U3OOUJkPLmbuQCcyv
lbajwfn9UzH65/KIT/G0JR9DWdaYyV9914wKqyeCwadxJTHxg4hWA9j+k8rK6kOo4Eao5aJ/9fbW
1oGMsEHh5zOLsIj68kl/jv2Izx8UvgRwpjaMGKhZkvS21cP5eB4TYr8MDJp/msAlRJqfvnE0+fL0
IVlTnVo8tJyHMb7nD8QJDUmicssUMFKB/mpYLL1um7MqbZ5C40EpxMUk1hDzZCt3DMjMNeL37Q69
Zuf8zlBkJKrw0OQYkDieRpz/7VD6EPfCIFwc61WIUriUC8tVmmNdnk6qIjouw7Ij0paSXRPmYmbZ
xfO0HXhHqKAq9PdvAfqPwir4T0Np9HK9vsfdAiLW2m45+U1BZhqcT2mnyFKBox8N1hyOrxCozVAl
Ia6IelEhRrAhclydKOW8dyCtQ8//TIIXP7fRVF89pIu6K8YjP4SfB5zEMEd1UvGYXHe/pxc44bt7
OqcDWFeeB4zDycl4IAkP3qnWlqvcKcOGIsTD/QD3XYuZw3ymbvFgWB/wiiVdbDRyZcp1Id9tVju5
4lNaKTv3+Vh6ArQSZL8ChL2RwqqpucuXSwW7HOjSx8Ty4Rb7zCVMGyx6RP1gO/GkT7KRlwAhW7Ty
e+zUCp70xoDUclCZs5tivVhFj0pKPLxJWnxhDmsb1sTkXM4tYinf03Cy7zFpbWUxjhghPmgd0w4F
tCXy7IddfwSj4cuz6y0LnW0tiWQZKKJdhW7BoWx01TXSkiMxiGyFgPCbOAZAhfV9Xmr/ta861Zv6
1Brs+O6hb397fuwZhjCbubRkByc/IbxR+/0/XoLUik50GNqdzOM+PaDCW0WPmXzJ/SdLDzU7NVCZ
DhZFxWSHqGhxcyohUMLmYz7AX2TaQ7zBlmsvUFIjTdxNb80SH7tGsdKrYhkhSUFdJZ2YP31jY/2m
6aY+ZOSS/CZEB5CyTTyM5h30LLvdZsPEPmC1Km2iJ6zF+l/eMCkjThndUlXIVNQyo0s1sw18VACp
wMGQaVIIq5mIyY71ShiO5IOH/nyVs95VhyDBbZ0LS1MzkgmNbjA91SdmjGXD7yZlull+X6qiAvTm
A9p4mu8ZzB5iOhi0usc2+etiS2+zE2Q04xsf7yZuRpy6yeymtvEQoUZUxdRQaygofyb5oBV2bW2r
gX1PbC+atIXm1OWCr5Ildy7V6ncLIuHYQW+CdfASsLSEq4DzFALVzZJzcg8kerWNMoRZuxodJGLo
biraJa59QUart0SRja/trc9YlkHUFgN0b6cYXZoNY2z4WsmzCrnWUuTlILgm5ifh3YInyEiAi/NN
fKn8mvlfpvowNnMVFQFI5LEgXvLbWDz4nu+E7prdT2ncMXTIGMFL/o6e8GP4TiqPO7keUBmgUGKy
LSi/W0lrBrKXTvr47hkH3UXsGaJvSR7jdhWdhBOAU0qMjnZQgUxMxmqsYjxey2fDYuS1yS866RhD
wrJRsWEs3t0IxgRuEC4NhrM9hRAb8lBYjzpKSOJQ46QtxK1G4J/kdJsVoYN8bGKmvdCcgfEaFIev
tHbqS0tWP5hR/Uzv18epT/fUcUc3vcHGZPqwZ1zdyJR/huLQivdet2P3W9kYE7IMdvRguWnSrcAn
oJhER7O4ap/zQiCLhAMjIbnq2gBux3zUC9fWLqSpASsEOVjh1wGDDdfcN1vjVPs9yObSyI+VEOhm
QtKm44QZzSlUqWQYoRebDnxE5qjfDmbivezil4O+Zb7RKsKchinl4W24hGshfWvGvlYtAj1jZfBD
Ovw9UJ74CdUxdi3cVC80hagL4bRlMcqcp4RU/6r7f8l7Ms0hHCD/qTgQKazuBo3IeAZecDqeuZrC
urcCAO84lYFsyjJZXjRJ3gDIoyBhSsqYxVVOtEXkMnrlC0fG1l+N14PdTTek+N8VOeXDGEoF7sTa
S7N4z9judxRlxR4tI3w3s5s0U5HpiI84ZB/xc2qy1UP33g0+CtzykTryCO8YjOvKs+a/UlOWAqJL
IFX92aAUxeFFZm7PFPYG3ZJ5jfE5qIPKCUG2bNGtHqYcMdZzJh2rxjL0R153IK99upGiRBw6InZz
98C4YRdaf+l9S94Xenw/3mANDhO4z6Y5iCYcwa0+VNIQfWSr6cnShlguY6bSQdfTRHUIfsmzYtyC
bjfK0LLUiXc+9ZBuT+lPgoeHWa2tiEzvvrurqCKn11b0kdSdpyla7ikCj48cB+CCCbwB04767N4b
WSRWXzNTIM3uKZTRmGHFek5Od0AMULAkI4aTL+1tqLST7rc3rmN4YeMoNmJAes6xwK6B5HZ+i3iP
rdnn1A60z8dMbuw3eeq6+UTKhFaG2/SuyG2b0ZcaHVUpFTswHq0rNPSyCKQXoY1dH7wdScarxawK
ZKvsLxjqz7cOc9rStYzpgWVnC23TH2ZeUjR6oUrn/PVKCj1tC2eqSbUz7IDpRKczlELnWJqPbsp8
NENmOLMi0kfJPj6lZ9PU9bpBk96rmeEKxbe3d7AdGnng9umJFs0D2wTxE7SFHzenXlFiiT7yy2Mb
It5HDWnkGkWtRdutnGtXFPeq+pm0qawb0e3/UojCn5m+bFIydi5JRms7OVzGHVVjldChFbYdeN7h
ZcCVXuTVhmEw5UGSHg2b5KRseUiOFsQ2MP52wUI1nD3IWyqRIkhXDvUxrel1p/iN0F8c7S7QYFdW
N7UDcc9xddlOQOmIxhrZnjlNPrzi8A5kQ/QXfHSkGPDX0r71qkWSDKDSZReEujHbjDHqXZ7yn82p
APOl5DT6oN/O6bcp2a8bX2uNXkm9NcMXH/vZxwjKgFvo0GIrF5mMOxRnXmwYQMs4XiD76iVEARCB
ncgsseRMRxyymVtHqupcnvxVVX3VVusbEt/L31BdSKbtlFtwtQ9EfEpsE96aENFDRTZoAzrbkPXL
6H8AsGRJXmsu0mTx9e4D4qcJlxQkHFESR14cAjguND+f7YqVijkg6zGNTyPeGhjkL8Ei27KapvMF
omEq26EFJ6766+yJzfbicTe0vxDAzdnqh8YsgCQVsrVYsjd9YxmU+sY6ijVmKMsuOurXWq7VkYQB
QwKkYeQcIzXhf9mlTG0ibUkZ1FoLgs1SQ2yxI3pWmU4pErNxZtCXIa1ssA1x7lkFSVwvDRz4R0K6
w2XgEINxarWBB7Jq+JkhCRDWXjVltZzXv7m6ChZERXJZxA7JLVb4xH4+tJBw51nExPYE2e3YsI7D
uYD20Eu6HwiPORHnFjd/STdBOYA04g18+QkLKLPfkdQ65b7zC314wa033E5q6H0mhlJDWdVT0aE6
+wyvq+/X9t/bPoStlkmmDYDvJtHPqs5/7D9YlajUSFpoyW0DmBTJ9+SiA99Om20m+BalIELh47dr
UFeAbH7GBPz82g6bNTM7GTxO1LkZwfEqt1KGSUA7ZM6ZxK/9A2JGrKIddlxg5occIarh6xAjzlol
n/uB+TWAU9UMOo4cbyjwx0POcMXgAFtOjx4De+1A1ymzshLznDhuSy1i+Ni5qzY4aaK4MrfAHl57
h0QBKARxDZkwX8613/t1mptzA3l3UY9xvgUyb29Wp60HZRB/j8EfTgif/YLenhxzkh7odh+6vxmg
FiUX3blAphWsFnt1V5nDjLtp8fqFjj1mPgA2lJw3dP/20naKQojuC/aqJm8uYTz0Gz/9O5R339nN
n+pu2FxJlE9TjLYFD1xUIsP+gZreGrzeXQaENw5enaAWnUyF+rkdjOLflwRe4Lfon1rSURGub8EB
N6lAS6f4RMjiYoQgCo1t1I1hX1s5rLXbhfK3dnZtL0+gtL75vUzW7rlJqgO4ibeD/b4drsa1Lt5G
NDpoLWTbt/7uix5PtuAeLqRzP7usr1L8XkMnU7P3Zvxdf8Ki7EaYt3G2UltWuDX8GD9bdsDdufwz
3oy3IiIlpl/VKdekyidRnK9BJ4+ckNAaI3vkJt/eOKkfy1KRwcv9nrtOFpATgFHTP3qdV5Qgvsfh
4+y4sDcWrDeP2qZ2hgE92+Dn/fYkfQJtY4+sZd7oZ5wE968qStO1Tdd0h8dseUzqyJYQDvD1Q+iD
5OfMAdeHRtr10MvJXZtWgQyBydGtrgXFgS4A/qtolNNfzDPEOMFlTBnW+zknyOpM7ksAKaSHE/lw
AuRmcwAPMV+e3Tz4Whe68qRsko8atu0C2iuJYbGQyRASnW23xQSXFm15oGoohJFe546SOhj7CBe4
oAsH/0un2zKEosWemFoPBTZ8KyloYdY+msZK5ABtOjYxZqHpVPETqPYz6sSjuxkP85QSxhV5BC2F
hHefA9tfglRQKo8UIzhWcQZ4cWmR7s3XNjV3YoGZP5iog/uRqvERmUOBk6aAVv+tIp9aj89E1k/h
akoANh1xqX3DXAC52SvhzSNnII5Ae2a149yzKVaQrQ0RKoHfmueTgkPvop2d+7ys3a3rfqQPvoNB
SNazXmvxbN+Mhc9MYfVU3sIQQnZiQbtehDwq3QjvsDPrwSje6TniNbkpCzAv7zPVthrV3UeRJcry
JE8XYLUcQQkTI1FbItex9egVMuy8SDt17Usfo+J13mu+2WksC2XIkuwbjmnFl3pH+qmdgYWxo4Na
l0d1NqnZjQ3o9Tlt21PvfXXFt4ZBtoUrK13y2r4nBWBB3rsvH0tk1amTkzUqzIWwS7HH+pwkNZQr
MMzPmxVC3s9hiS0X+puBTxM+BcGJfU4mi0V+wOM2XoMYLIgcdaHP49dfOvfC2bGYOXWJV38axJ8c
wIcWqXL+q1Mb/Cyc7SHD1Cquh7c/YJgzd6X4P/UHbTGB+SI0r+nJWaHul12SgIuuRmXDrHrr3lGY
/f9qnKMQ3hv420WROtYXI529k3DybNTDe+vaMEcCzPges9TsUUlxGyw/q2UsKjM5sBl46SYBYARs
5kWELvha9NUTIbxdzFjIhjYvG69i9aNRR52679tTgXolyID8dT3zhl+o1dFb9JktTmb+KxZFtLVR
KhiellWkC5dfO2EOyjzteYMBAFkEszNtPUeGZdwWH7oAoK3+pJJklEUzUnGQVkjjGl311ktY57GU
Typo8ropQk7uuJYz9A35R3r8Paj5OmFRtbxJdqEk+pI5wHXzHzuN+/Zloy2jlKe1wa3Ok34bIqzc
OjzX2X1g8E/zPRrW6fk/5tpeXRu9o4Awvc47zQAd3Ntvq+Q6s/JViV/WYRq8TPBAEc9i7eyW1Z97
vmTIHvfDKeNhPz9wqRGabW/6PO9BQ0w1DmI5bXLGAT799eAVMQ/kNRleYGuVwUDQlcResc9mbAMc
V5D1o3LiBq66alQNHXk9IAUXs33exYfgwUEkR596wFytGrLAgxPTCxGtougGF8iaLmkkznJX2sCb
TYmOjFN9nwNQVpB46v/KACCW3Czv3T+rO17MtIgDBFKiR7zzW06S0EGld6/BP3sIG3hL9zUQI+0J
T6S8+voVi92/zQkM/LoRP7eWT1fY9PdvGM2bHXmKuT4XvkMRMoEBfT8IxskPc6XcM+qnCWMoBa7k
HQ2ORW9Nfd/3GIy+XJodDZTfWtG4jH+QBPnppKbZ8IzsmRYw4rAd+sfqwpLFbd5BQ0PDzWzGn1hd
r0leqxO2TGbwDNTutBmAFN6OO/7eTQYMC6r1u2BuLd+dDxJqrz/Mr1dhSnAm0YRlhpJz1KGF+7Mt
JpxoCfZvF4UiNOcFJW051zjOcCnk05FcsGLWyxMb+5i2JOyZqtTHHEvS2OoKrQjK0yICkSCOAeIB
aUzTx1fnDnynviddz7XuOf72Je122SptLV8dlOrKzeR1jSGdhp6AHUwWu8w1op3td2+sUB6CgGAw
CclBCHclRy+TaoOMYBqDwh04OVy4fVRLkCuaEey+clmT5tn1pA03Jug5EyFsvN3Z9fMjWpH4rr42
3jjfDXBnM6TdcJQaqTuw8eqSLm4+ZoOwb7sodwc1BNT+7VQCqvCD9hoW8CLhRlxVhN/KiAONSsqT
cpuda/u1kNP4qeRtWhijYg8i7Ej/OBLCO/5/ET9+6dGvraen8M6YwOWUT4PyH1p6z9za8eQECGSh
fY/zGBAWbfT5FdqIgq3GNrp7WwAP/Nd2y+Q47pE/q/KwLUfsU0H5ZAuR4R4T3ig6MgsX++0baB3H
oWfBsDSwbSN6blNpV92ULRQx0EKPrqjAUv6R08kX922bAdU/hbgqNamhUEp9mOh8ZYAjXUwurCEh
OluJOqpm47rwaVRGW0fhwD6n7qWycM0ktEYJd8nnjoXgOqBZQZo4KCGTwSR86iHKCz+iwy03wKbb
KUrHA1ldmHg+pQ3FNHhJZzePRCXRI1fDvwVGSEUTkgXXsB0w9yAom7UgMKh90ZFVz5AfJS8fIB7V
POIdeQMTHmUYuxvgZORqyXERZsBXgDuQ0l4kz6y3fgVd4UoYyCdSaJGC87p7+ZsXukas28S38u+C
TYnmur4pGSGPdpByR0wMoFRCdR2ZJJwVMnLc8FRA0m8mXZB5AMH3hg/YQ1AYRrAw1IxAPAvl+CtE
1q0DqMqJbbelSVYFKaemCBkxmf/4iN/Hdc4WP4nLbLRtguJQiXl+2p7oC2E92qSOu4CjX4me7Uop
f3Qi7nCxerjw5J98W+AbFjoYXr5hCk/16dWXxDUF692B8ZkPDeBhqjV8kD29gG2121XphLbmMhDd
YozWJIMvZ81UU81fA0/6iJPGTi2ZF5+/farnf8egnegp5ZABk7OajJjl/qJ+LKZwDY5DJ/vGONU+
SOA+rIfTRrLz4eXnxrlRy6UFBpwjpmFClXw+KzKSVQZEluEbuY07CoAlsfSUzCx1tC3bzeHlm5HG
vjDhkYH2Wq8fun+Fc1zB9PM1j0oaKRNO6m0puUukWiIEvkWTaOqFXkg/btUfIeLLFU04COM0z3QX
FH/+66B3HNJGcu8h5GHvtxm7nPowOVWqyhhq84Pxs1l8CFKgmSQ2XqIIYZSjovUgZo5CzKlE8m76
ueipjV5UrbQ5G2KLUhmAC2a6qxbpAAdlTeAS5dtk9FALnV9CZI8S8vSGTmGGHGzLwi6uZ90s1rBl
zfZo6AbSNXdWgWcHgVZ9kkiqpI6agUFrBX00VUu/lX3hQeRjXJqa47QpE4brZafpXCnaKk4rr//0
GZ0HOYb4LPc0de4kvfaNzgHzkNh/w2HD2sGOPyO2Qt03qa3iu/R+A78vf/lvnOSgc1z19GD0iuw1
PsEnmr1Ne7fGhFFHyhLATB/DzjhDZ57gVMh7BB8WBQYe0tK2ABR8B4O8dc8DU8ke2Fc6GwtRGQIk
P6u3l47jPjnUaJSOaX0ZHuNGeaBQOL0jtiXvZQ1G3OFMe1FezIeWaUzltlAQKkxaJQYuZ1qatnwn
1aqe/ODjqgQ9cXpBslk3e8Sk+8N7eBCVuDdOZ7VmFsdmfGldk7hzkJl3WMvHaDlu7e1YKRRmQybX
CCmJSWxap5MxHXZldAu7tYASPK2qx9qU5SzJPOUNzPYS4LgHra2onkOk3WomOHdNW7Wuy1BPLp/b
uIEEM6vLl0ET0/4EtfjJcloieR72fteBc5GDiqNDW1FRayMnHSdfxoSg0ie8C5KctZb2VCv+K/44
7rFdZdLHy8KUv0APZ4zQKh65cOhgB8t21uGfIU8gFgU1NgOVLg9dt5+d5S2JRSteFy6QsXRlcTYi
SBOBxXcp7dzxLW/SnoFkO4PWgB/025X1cMDB8spAuDklYFrTZy/wt0gXeYP1L6eC/Hx+Y42m1QFD
uqtT4Kh2m56y/Y5/6a+f9vmUg9s0PnUAGblYzPjQU0O9ydJvp50ZBbM/eaPrbiWryormt3udHxyi
CDRlSdWaGK89zdRICQXmyCXwuNsLfy0WCr8T5i5LPJOcAlOtXSYQ04IdjWmaRdN+lqJTvpARtRdB
1C6LRcnOmL2EMN4I+q8xdc1R00uj24t5Ibb7W+kccYZbQf1+gCcMEWwBfDaeVk94+riMAm4vMWYW
bE1jjRP6g8QSOs9rcuzxn+PzF40N117thffaEJuczoBJaS6R/+o3/S3ckUO31noMdjTEWnVOHLAS
bkHlZvDBG0g70CXdggX2IKRK/kKgxfbwP05eJLIggNRgYdtSE/G6QOV/wYufIliN60Fr/Q+Nu9Ta
B7AQYAxboJCEYJqLj9s5/tDKnTBIZqTBXCSxLil5IELxgi5c1G105Wb0c7B9VrFauLMZlYh3hGdt
RcE7s1C7i0KOznre4FsniQc4lBCYPt+7g+yfLH5NxfpHLkN6W8+e6jBgdSNOZ8HuJZ56qO9ADOwQ
nLGBRCnnq69EV9PjqBFlpcuAqS5N3VOws7RqhmWbxPivbWUhnCBeZoGYHoAWzRLmmobPCg3Zkq80
VzGi1T8x4/Pu5Htut2O0Fmz2tW4wZtrtFWTiYN2Clrws43+9bxvw9G/c8tzeXjnoslzkqHKmvr7U
Q3I8dxJdz9wLNzBinU+xWs+D2xqmhlMjU1nIx9lhM8QZneTHmijE/epV42RaklEUNVa7zQi6kSE/
1Yehq7mfvbETyFfG9/Vyj6sVWZ9M10/3Aih6/rqokATml7yasaJnRlmF9WXm3wg4jgrfh9Gbxtn5
Y/NwKCSTqdAQT+gr1Oy6ZlOCcfRKGPHWZhtL2CGlQugFLoFPOj61/pHOqZ5Ka2ACY8UDSorzsssP
HNYVL80Gz6M+wYTWWZJW57Bfm1fh4j+pUohYtMgm0faFmaBtDVa30oEBSRBE0oHq2KUPz0mi5o66
KuqizWSvo+nAvsMpOk32BPxjseGo3mNq0VKNbDIEex152Cef1TxU4aFOdpHO5X+xDN/NBPS8Mjqn
7XthuRkbsjdOA5fyDyN3EVyW5kSXvXeT/lG9sPyUQgq182OSWPK/fgxD0CIlBNWXM9pwVE5n+2lm
SsfvqZnSGj+7A2rctDhKPGj8u6xgkn8g8Ro0DXT6f8q/TCcghCbUWpqTFo6s94lLZc81ss8rTZOg
pysythPBk6spQwQhssPqCouNih3RVJrPhPpRCo08o5NQAhioY1e9nvhbSak9If+eRQhZN8Q0I9JA
pjwuJYf/c16bTSZk8/xC6YgCGT9bjsdymOgR7/CPJWMumY1ObWJdLjT1KKxxYkxu7ZkKOHDUH2qr
Dyt2nVQnpx06mtVndNNik8eui0nbaP160XgiVBa2SHnqTzEAGgeC+7Ryt5NvrlpvlpbOHNSrVH3P
ice+8v5M1Nef/IEfB6I5sNRF/DRn3VVGBJj3tRiF1G6DwnDLg0IDJqcDyska/GVNQCmb914N1+4R
0tVPLuBYJVYb7niRTd5kAw9/nWud+dUvv/Hxt+tGIPkajwM3vtesqrCzYSwCKvdqRmzvhi2EHquU
rllOkBYEXaHy2e7IBhwr/DF1PpiZB5951vauH/hfghvA3IJProhbFxohwp6mlDcOMIcBjC5sNa+8
JbN24/R3ZIbM3chbx9Rtf2AG4388F6KKcofCBxHZePNTDEd1y9FIi1Ib98o2c4krKKxNBw+ql09M
c9HjQgh8htcrGGdocrlfwDAj6OxT2/VHvdWLPTNMrTcaIwHd+175vVNJ08AdfI3SpVhFvWkTQ8Ag
JMg7z9VJzT6l4I5WyHX2xTjEJu30hCKzkablzq9VzQH5qngX94gGQnIrvMO5VMXftRx4aBvHCqVi
7IavBoG4HNPnA9Hqf3ScImpll7++5j/8ampEFmj6Lkg+Jh38M/KbNmRQImYlA8thEuu1u8zR94BT
M3tpzMy9Gh6XSNowp0QlYN2DETTXR2hXbV6OYu19ByHdyiPa6+z9qYusfSBP3qAsqRghQYAFqlX2
y8R7yfz/Q4FJoGJkA+dd6rlylRsbELDPUDXrEXwFYSZc8hRIaK7qWp824j2DAxBkt50fnSXFGOTr
Zp2X8H9a3k73K5fld6CbBNX+XmErnjgA/xy19C4fglDiul4kysqOa6YHp5DQX8Q8mnipVqFoawRu
Px/XV7vEB3B4t2tBQURmO6I9DBWdsFZZrOY5VUflLgWTjyScawlP5RHdVhhHV8KzTlrKAJxzzUlK
I/y2dzmgZWz/XfyzEUn+kbkOhCTiH6FRGAtq/zTzblv1m0GUKWxnC91YGxJCvuaD39aSclnyZGY9
E/Xq3lnBjLio4xbZwGsUTC8BJ4kSKfdaZLKKZeXCaR/UnaLbKYrdaGBz6kU/HANXpD4r4TGvTedF
w5olvB5UD1aXQDMsgAwXl9dzk0FroSbSsLeJ+PGEx8ciA9yS924tan/ux7Je4EKNp1j0fuBW7PaP
76pJ0wBJX3YmYsVqbgpGE2lA/5xvSpCpAhLmx7b3o/uHntISYv0CEKF5+4E1MEQ4x1IhZP+INbRA
4JyEYAlvQAL/6vFUjo63ztB64du10VarPIQj6/pVhhbRX2eH/Ye7fl9pxuE/rKMPx+j1lb/fJupk
E54trtRU7AGJSOYv6/5v3E5LGqtR6Zcq8bjvKGViwv2smsmmGmsXx4kvoTRafXOgfCIAIvPtvkG6
5U3PpObb45fDCEPliBL3gNbOy4kP4yiInKJdmzrmgw/GWFKv779TWR40/58IiNwy8EAY9M/uLRIf
cT4GsbV03KYBdWlCWm7Ne9qV6bqLjpcESjg47ryJ7CpJw66kh45apn9q8DjKm07F/LqEJWE5AqHk
FDpuBXHbf8W6AHFeKxDpcDEZyPuSTm0pPhkrg86AaPsyMM9o7adzuF6+GQw9yAjorAMZ8zpQ1k78
CArvHv859DIBK67heIoCOnLAdf5qiufpOywWX0l8MZ64mJF12AWu/xB+OchdYl9uoLDyTchtPJN3
wtzPv2cT7fy1uEyhh3PpbqPvrhl6kJp+YtTK1dB5DMj3vsE5Cut96fgrZy//cTVUe1XH8JujrZ0u
TOIpsChb29lWBMfSNsx7ELGxiy4gTCaraXU437qJLHyULv+8KLR5c0pKz6+9nrbg1/x4rv5yy39e
tLryeXyJgYdgrUeA1ElqM4cob6Qg8/KfH1Ahn6cnVNh6vVQEhSGn/1HiEQnHYS/oLyeYIF+Coljh
MxiBeH+u7Q/EQrKwb9z/Ru44QuQZR1Gz4CyRwAjjA3cGu3C6+8cLfpkALyHCyh1JIY3LuU7ViopB
GQ6G/97afX+tcwPNodd+Z9LFtk+0cNGRzxa1aAtRp7BkAbxlnef7I3T+wm2f2mnkEIdWUkGAnMEu
2V6S/GkRX8Xgs8GcsLef3Iuc531jL6DK0UrU+SfRWqQLIPE2E/tf6idEj3+HsZod30qqEqf4UWXr
oTskCmjsRCNKhw9c9LgL/e3fh58vFHI7KbIrlXZEtjzd6GNs/4ead2QHv60USNjTQ5+LxBlPF85Q
qj1UiohHPlQQ2z/SIDLf2LZddGM3H4HhSaSCL59Cetd66MX8NhJol/TDxdwApKqBOhW/n7AgG3bC
L3QjZqY9cBCfW1KXIxessFA1+eiq05AEENms3keAEGhSNUOXTrn9ovxtQrl+pNidl5H9kMfZ+gf1
oKM166lh+M3EHgrpJk8DtC0bZgVog/3mUQ8Zicnv7rrGmh6LERBTiEWva2bIpMlG4wcddBMJf4y3
rxcd2plX0hLGnKuFiXTAeYieuT6VV7RKvpWgSTYD+Bp7g9Dyvg8dcozoLQ9ImFnKOOFwoVPesuAL
AGZ5LKc4TpV8CP+MA2G8tX0GqcrSBps26RVSACLHHqSogTQkOdLM2r5L0DeF3+UzhwqnblNZUm/Y
GTl5sAZSaBoZPrMGIUKpT7jogtauK0qkkaAUjPMRyVRK9ekONBgbYfOhyS3n5mZSiUKZ40OXVSWE
NgLKjn/lLUa06XTHJx6mifTvTWw43/EdA4Z30n1UWB4UueNBIaGGFVifnRktfa51GPJqamgwTuFw
MKyRuEGQnypWk8KInmMBevCtDuaCpudLPeckaoUmuhPfxfdimRSuvu13kd+RYeN3tautIQeZB+Dy
RRrSFzr70ECKo2P0yXOLfdZyhk+d6TWfbx4Py5+NpR2whiuY3Eht/3lPg0Db2NwKRMlsIvZGy2Jq
iqP7NPuwtywBuSDgwWS+pwD2+l2Sy2o4/KyztyApnZZMpCIThtEZUyLGPGFfNrWJlUVp8zD9Fd9f
rCdalXopn+VJSDwJ09T/tnjWyBv3S/KHZzOpzoEWodTL2k50eTYDYETBDQBypnOM/8qNIgMPrXoI
INYtvEBzLzMW+mXA2+D7vVbrRBbNeXplTAyS7DO3TohBFnLt22/cyPM26T1gX+M1xa8qw7KwwCV1
H/mY9eHh57knXY+ADf5R8l4kqgqyLlWfC/YJpkgk03ZX3UtEQ3/XY+FcIISIZDU/mD/GigS/fSag
we8t8NmzLeGKAYkUHkQirzxT+MjiI5YolvBRuxUTB4Oz8Eaf9ZdEReVUNibVuU2Dw2HkUfB1g4fb
CdRDa+bt+OvjKCv5YSMr5ZJa1Q8ug7qB9WjENXiKY9VL5UpUBziwsn4Vku7kBrEgW711kxR8xDjt
yjjqS5PaAlWFQ5/PruzWd6O88ILqgPSZpnGKPNZRE5f5oz80umDPVN2nxln6thmpFprmGah8lgjg
skjYPs4GZXrp4mM7Dm5ooUWBW+1AaES5c8MWiYhryTF5ryeHedt8FIFsEAHo0dhHufe+1NVtYRZL
K+nQUWX1u+JslVicnft6Fr7KDA73bifEb9S8AhraoWW+/4ZE81ibIxxqyYVEnClzACuVI3q7PRnV
Mp4+VthCQ9+zSxtmMTmouIc6czcaeRC8dkh40bGQi0lkNuo8LHzISx9BVVaiOiXbPnUN84d325eR
tUbXsav1indl4wGkNkJ7Zk1G5vX7layiiwzfK/LVRuLYaHHkgMx1kQYKBaoA33+vfql1jDzAPE0L
/KQmht0avRRvWl7/69i/Pc8d1QopnMdBLe1EDpRU8hMlnzjcuHq5AX+Im1lTy0qoi36TWmO4qXC1
toFb8Qk0GfIz+OH+pIZVdX2LRtXXntnCPOXSusIZ1wKEpoJr71c9SSih62RVTevzugzIpdrLHRju
oakXcCJTXqMDcEiK+zBH2Rd2amhxJnYqH0XDh2amke3BvDPba0EypZJ/v3Z6TvRhUAjxvlg5P1+U
9VzGSSm24baeMTKZ/ovIVg2iorwIy8/758zPVJM6HlInGg9Wb0NiIsoOjUkPe/4qZ1+8Bxm1ERBO
AEklKEdvJ+/jH++1B+bOg0Z7YiJ/k9n0OmivUFIgvTCcW0DGX1MTwhDHtMppt3cp/8SbyLFIcybo
vxJnEo1yJSRJHohWfgBHZgmwdRn1rqoMYverTxz3KbEqz51r9qMU6UqDLAyhzu/jcW03M1jYrKtc
AQeqxiriTDARn10Ush4Unr8H+WhBPDdRhtyg9ZnQIPzWwpQ6+WcztmTtD4FAGizkykvSSIUOzqGz
0bcgZQ8FMZFopdamCdIAJ2a1j2cdrUkf/oSHfkY7u86vKZufbwl94J2pAOgge6VHRqcpHgDNgOyB
SxDZAgpBZkWRxBOTM+q/w19H+/lWNtlvcVM8QhFJPUybkrwifuatSt6uHl0rH/fYQI/KrbdfiMdo
YzcAqwPoakO/uSKT+QyEJAXzXUOlzGrmRWRqK4QcefL+NbFNwVi3N9FIy0cvdPHJZKcrKkbTR7+3
x1il1Okp67qgiOV8s9I5W+jgthoBTqJKKPQ2eDrYwwhdgUruzC6FhjDy0JDhV5eVtPlpApnXC7pv
1KwZtVmGC1MoeStawTlhug8uijYRPx7GGfBSkmeUP65xckMqDtvCTN4c4k5JMN2t/912b4bDYRzt
ScZJ8f4b/IcEoISFZUQR8F8l+rYw2DDYdg2Lvb7LRnYYW+Ln4PhGAr+VRXYLWCGB/SfDZd24Uqup
SWTw8kEtJD1NYMsnSa6MgX9VVwytTyvG6RmSw6znQfy8ndAeB/rdMGicNnSUQd4Gt2/2ctFjB7hD
dpZzDx5+K9ddVpVkKNSlp8ihM1lxrxw56IbdwU92CUBw8uN4DLGfx+h8Upg0PAg1mb1Aw397HzMI
833eVPLFpPMRhVc+EWOEYaiptoKsU9PXiSz8NmXrqb8wMmW7EHDIhCX5dP+v7W0tVfza0xvswjZD
bzaYlhJNg6MksMfi1+CSUOCC6JsHkn65A1RxhWlQ4UvKvQ2RU+ViFmjWxnZpktqD9BsHfoC3mSME
78gQJCtrtGcU+tfije7CC6EcAX6xB2B2tutHbD++DgrhJFANYyr8wd7Ii4FDF4nROBw+bmZp9fu8
XF1708H9SOe8lb9L4vgWp15tjPx4jHCjqqHuWgp7PZhJ3gmnkBZ0YYFBjJ/KzYhY6iezWNv37r0e
Leic13lhYxw1eRI2eMDQdEGfGugIcUEE4zsJeJO/dfFv2/0B246G2B2wKOSEJZQT+yeX43uR2Kce
J7NHuS5I0bf5vRIkKpod1p/PSZvH32zcW57JbI/OFZho/hq1aNzcSQbFqiW1Nkb29KpeLaQueneH
GxmiuXxpoUDbJwrU+63e0yqcilGVb+moIX9pqspwYONynUOiMio0SKsESNuZSLrosIWqI//8yv9n
6GYbVeuo6AVifAuhO/FGHNa7sA+EzopmwDMEJSYnuv895W9DTWosltLD3i/cudoZPHAqIfrICz5Y
jdwhUNLF1VZ4q3BORzunQyt91IybI0wm0kmVRCvXGNww6WNQF9ZlLe1Q4m3pNZz22rInnSRj822z
YVTK+UiRP+LfTpU6jaRa5jqRERejH4aqR4fWzSfKIpuInPJiD/nwYAgWOV4jC/6k285zRZb6aulp
BolTo8vV/WU29dX1qUHgJ8JKfoxUm/ksOuXnI5Mnqp3fr5cnN+C3aDRG9Pak4GS8QtA1ORYMXRMd
sGyujPDkL4ZSawfCMAoS0mVPIyqjAkD5bsF0aLeh19UCJDtmcVaLvBxptzo9WRuIy+dTs7HcjLpr
3c/PKh9wYsvVXy83m/s8cGu4JrUuQiXRTZkWMB3IabC/1cVr3FdXl4m5MODkd/OikVFzeLOY/O75
11VhVaBGsqFUsOa7ccJ/L5ubR2ktS60HwrI7TvgXTB2UYleK4PNFDJnYm7sGfBmyUFii9FfqvruO
qiK6iGJbMWXekQueeEMLbSXtxDd3vE3FKR/rWRxB+DT/sfAiq+grtx7vzOzLWZW5k6bi8Qg7PoDj
Kd2ngadphto+U1cWEDkaiUbQs2XIQhr1LIeceTHZrsPpwUoqBTKXXRWL2t+Jz5z3TTQyPbqjgYPO
vKLZi7CM7w32ZyarO4cFF3xSejH0wYLviYto2eZEVyNSMSm6qs0a0I6voX7oRLSS/QJ3TmFYUoqZ
ksBDWg20WEyvnhFftnc1jf5dRqgkWBd9X/tomTJcg41PYNv+2aCwK8OXp8jjf6FsFTO9d/ieoljV
51UQDCSxwsddvYBv4BHnjSxOPfOSVeRMC6Z/N6gBZP2Fm7/SJVt2On3R43ZYpp86Q6iKA6vTwCGg
kjYVQ8Mj2rKAmNkmWIaXTegm4zv7N/+sSRn8JTJqM3veV6uHWTptrwcT4fXrMRu6KuVP1JS9KvOT
K9JpjER5MczkTo5rFU6M/4cMe2EtHhkWf2BUxJlX/NH2uee3qvzHprF7Qxm22owQF3aSDPuYn8t/
n7lYLghBk/AiPt/gL5o7t9mYcR7rXuZdK1qf41nydi5N7hL29h0/N5qwQU50Y3ER73GZTZOtSVlE
PTB23C4EI/d6vYrkgo2QhnWA55nDn2A5cptSCqLzZ6JRUR6Oem4VlZkhpz+5o8Lw0cjs1uYccsTf
5R7WJO+9uS0o31PEJKFUn0UtSl79Rg0vAeQ+mBxmOlfLCLParCpMvzjMZSQL0hawO/cheoFAqBLq
+K+iBUYtnZ+7RLoYH51K17+jTEVRuM87QQaPBKcnOCmSRi04Atwlzz53bVhxHxolyaaxggv6CiYg
PM+8ByoAYP4yEKjRYqe3dFl51e+jeokR6UVVqvKGQ6mhA1Rmc2AO8WGcdbaXGr/n9krhZkSmT16N
JEwrw9AvRUHEnCK6vtbqF6iT+cZ9dOOVWbvxWY2kETNPHEI83r+Sb6KzrKpRaX8CkUNygSJgWaGj
4ZrVRnMLgCFgPJwDKhhz847empHaZY7qjLiuqY5wIzSkqwx0l8ke+wHrbCi0Thymyp3OR1z6NPlc
BtSGKrXYbrDsFcI/ZjuOKpVBWQTGp+DiOk1eWQ4s7UEUr6u6J5RyV7iIqW78kAjfHefQdHwbN8Tv
aQu4BURoAPHx6KW72EII1w+mk78da67lmYPuWrBtj/qoVhnnims0xAyNNGcTzbdekVQRgms2wKq/
qJWA2nuqh9p/dWwM9VIDGIv8xu6zX/+dvMeghIKDB53DjmLBElxiwsA2ISMwCQiBPuZiL6eTf1Ib
HOC2LQLCkXgEXLofucrLt/wzt1w/1qTZEdhRhh/zlPmhwjUAn3xejYITWz8OoBSFmCHBxY/rb5ae
62+MRno/I1WCgW5fBJ3DG6A3bhQcoAy6yf60HwHgNvN4MDmZsN0QjNVu9loqfOUYTWJpPoLgeHyA
oZ4BNF5Bfbz2Yy49isFRGneoQ8kVgypolCrdxrgxb6xtyGLx5mfOwbdQgQerSnHyFaFB5LCusNxZ
fGxT28wi+yJpPOwZ5iu9KhmEouJJeS+t9oRBULxTHAXlJEltFuS6lw2R3Tiyux5iSTARZmqQm4fK
PlIwoTnm50XL0UD3vYPV2NK0Ayn2e4Tm8F2ALOB6OAn+7T8v7JE10DnbnnUg1v3LQ1bl/sCYD6XS
GHSkN/PRzBC9sHrFboK2i+hJwBuH+iMLkn0FdpMildRpU83C9uuZzxgdtbMc2E9xk81Wq4+UQyNX
egKVLNjVYN/Wyabye4qbDgJSc4UKuJJVApTEyBPKvZvmM/k4zhxdYcNBSgml7mIBFoqtqRdeH/6B
rCSwJzqphwYOgzPwaNZfBNhDmaXrCGtHhLOv3hmQMTYYyqhnmF3flKP0NCkd/hT0Uy1ApiOkmqdI
6vJkh0/ymm5xyjey1wHYPGKSv8h4vUwbjNK/3EAxmOajJZfw9yXL/2EVgrphxGsXdnurnOY4RyWV
bEF2WC10X1cNrjtjDKcnjGexmQjgt6O5Lv2ej92mzlqDjNN79dBJfoOhhfYDMYh3uxcemKqP5RgI
El8r0BfwLOIoulgY4fQhTjAxJJrmkvht9pvCnTJT/SIguT6tCmPv+KJEpjmkMl2ujVnBgMfYI/8E
3FnY4Avy7pcsE7RO43fCOGrIFEgeo5wuixaOCRGDvWWH4pHXYG+pztWI7S8DMALrjuFC2JOSqbw5
IA2Nb+Tl/NVkjaxvud4LVwajszmv8VChSHfk601GCW+TkIl7H9+tLJ42Iu1oPqLQa3N+AEakaU6j
0uO3am1TcN5GEIRenzDbhpAHcoug4EckhEtz9Zc9oKYqItW+vwbsEf5Dxb+raCe0oM7nlh7NFAIy
8eMg6NNF8ZCrUZZJg9VQygh2ZEGUgMg+uNp0UH9m7CfeFnMyAqYoxNtkhsjOSXENB8T1nT/jXGDr
n/dz3ICp+DOJlzADoMEdmFGDSZpvQlU49Rtw5gWrhGFfQpyWiX2UdyO/aKernPfHv5dljy/JdsL7
LTJZFhbvuhwjj2L7P2Ih5sIIRT4B+aorNcPCEJvLKCuOs05/pF+IlPUo8MTksYRyfOgUT7hG0gT+
xCNK6Uj7ioRbVE05ETkQtQhNJFU6E4J4CzoXwy9IEQh6lxQXxLg4ek4lDuLQZQCoseAhIlbEAXfC
RnJ0/PMLjONJk9CP2rSaWb/R8SeRooFTitcc5MHifVIsaQNIIdsuzOygKplZhL0ixPp0WSoHB/VS
eddN2AEOg+jyZv4T7qjtNRQBwVguV1KAtNtiHD8zRM5GfMILa6jUyxuJQkuesMOg4KseRNPClVw2
VUG1l3pOBH/Y7psuZOA4pfDokweynxVsIQpTlDCnhojDU0H3Oa5L18NZI6zbQ8HKM4v69SpPMSiE
nE2tngnvpzZgVqFFG6IMFYPyuPrVqeOOM1H4tCe54dTza61r/8yR1/P1H7Rfl6v9MQA4j4J60Qqa
fXbeIRl5LUV0cKRrCu58wd9y4GvAgeOjJVj2NbI7h4TWOzcWoq3sCd5k6Cfsop9CQE470OHHuRTH
kx/XCzc8L/v2wBFWPrt8IRx1PsQMQBPJ8eQzUu7A2xA9vS2fIyJv708ag5sh6JgEQHZuuKYuBHO8
F+o6g3lN2L/RuSwn+qIfXXqprGexhUNs245XTWUzUqf9uWHvoPfi4sP2CzWDUSllCkDeWoux5BKp
y1ZOLfdeTzpFt+96Qu4X8v9EC4qMQBHeeuIhNUh4yJxOx2BbuUR3j28spoEtH6Rq6JSDHS2SiS0Q
xtkmjCiIknQ5wr/Kvpv7o0kftIq9o4v8IcQ1tzkIngRBo0qmbicE2+G7BD4GZwky1n8XTv1FrjDP
dOjftm5Mtg6XuCPegld/2fURjUONUqATOTS8pibgolFS83y9WPHLJREF2nK/4ECbtOgvV80thJVw
8NBeThOwxo0GolDoaQtcc8WtmHfyM+HQNP2WrMX7iB0L5mS1uG6cFz/vwjPYUE1Flgdu2nNSbRAM
2wDneliorQRALSgn9p47z0/sPjyPKNwhfA9P3PXeLx1waj0WCTC7nu5twiewx0OIZ5xdI0VzDBkT
3FqdMV/3G2oWC7soPjoUDwbDrDUG5cVHVkZuvXz4Kb9yJ5HGPiixLNg15mW90oX8xQNtfgU0rE3n
nprlVR7HSvKq43ZK+8gr+fIXM3t9PWy8oZCYwdAfaCMcqyhQGpSWRcBnZNYLYcJZuMoXgQytb4Oa
IssJGrMjYby9QxGwVWnxSOzHjpZYb5hgdLqKgWy1dvc5JCjZ90IMOkPwyMNqno4SmEhWwguQkUbX
0BWESMvVds0GSfS/eJ0T4F0G1E054AybQ4PM9fPeeOi1hgShhkphPqaAj/R6xHOndo/96pavloY0
VELBJM+HMiQ0VjyW8lRWw0Behmzpr6bIzbxXboqbkt3e3jxaAts33EZqrbfjGIdgyRF+0vWosIx6
2qQOGTHVxqKzDLXuLwXR10oOiaKKFfO6eJ7RAZYonfJuLq6NAAotR9MW17uRIEIMWxDlXzPw9DMB
CWt9ILjU8dlrjLfU9WXrNNvXfCZuEMSHkhOsmqB24dH2CIeaF3c4tFt+YrHJNOrXHXrYJmtvduQB
TzLAEvptQA9RsOmWlq9ZLWYKfuQk8r/qC4JZVHFIJ3FYsFfI47OwN76WrQGh8ZYHzY07J3xVgvDA
E4MC9GezMWjt2E43hgSK4zXQbhwhLk8j/OzFQnILKSOd61cGmyWBp4fIoRKGzlGcmiF9D+lirHpN
UOHjGGXAMqZTecSRQVb8rMVLhGxFnQAqMjhzdvSw5ieMhSljaFaUqArVZPiOd895bp8d1YNWDfW2
z2j+veM2pQM3iB37RympCc+hmOOOctoOzaW/Rw0fqj+9TyArS/fwd0JBi3TbAQmoPrlIFD2RDPpk
ixvQYGo8qYj3XqWwJUCX9a2yIyDj9LpAaYTFeizSeLYYZiinnC6iDIifzhqYtHzhTLgCW//kxBf7
1p+I2+rE6UwkMJT9xyRhX3cGppGyZyN3S8GlPc3GoFlmu8E0vYTpTn9P0qR+YYAoOS+zflaD/mv5
sE0LokOIxiBKqMnrppXQe0jSCDI0QWO3SruGNAkMMg6oEwYU6Uk+ZKMC/K1XPhU4os2jP8cGHZiu
et3JF5HftxZ3N6VBE8c0BFRkwXQUy9vFfQ49bhxlFiPrrDaubuFYPAJUMci+zEBr1Yt5YuEbHri/
gfAwKM5B81AwGWgfpA35T3JRQPQsSWjfnwHjdi6lPN6hLHoF6yrPXP9W+GX1QQnUDgwhieI9C+Cq
PS9/HJi7FsywXHpXiGKUD7Plsju+QEbPUqgaV4j2ro92F8kCDV0eD5QRsO0Lpc4KUorHYifMlQyE
cdbKUYpdOscRRJsxQ85iwFjoA+3oaqEgHysKl0w2/UzeU77D53rFIYBkBNFE0mWHRrFsZDzHIlAN
k/mpBcq8Ea2WbadA7tfQXGMzHthdnRMIpZ9JgR9Jj50CGsgMtdvthGPaeQZdRSAhPdgdkimInzVI
srUm67M1KtZlyM4/dzBrOt+iqm2Ym83rouuFu8LtYQAnmZkKH86fSxeydhAIK1ARaJASzkTkZpHG
JaWgkQxwoAfVTBYLIAuNjYx+Hp5d4qdj4EGeDqP2Ribp4UbPfTVP5OZaaPULarr+PVOPjiUVJFIS
fbrBigWRvlWD/SKBhIPUwLNCLCdtKQMkY4kJ9zYn9Pm1uHlTcUDnwKUVOiCDok9KT8FJ3yl3uh20
bvYcBbNp4mXNxowQGD/jjJ//SJDFwBtfsOQaBZIO4kx7ZbIQGxnUqsynfHyDFdaqS5txNCOIFlAB
JdC+JlwcKsS1Aq91Tng5qpVeseChsh/N0i/xtuDP2ttbbas9gdE/wluNwK2TZWpbDkaJr+j1VOB9
+Q5YhlaDUH+CczP8AWUQ+FHXs5p+ECSKaC9VmKRyDpRzbxOBaBUmpESmmSk2WRqbYy6VK6Q+MCDr
HRRFvfJxMUNF9ODJv7SfjBbbbnZvBlraHgXEAky73PnL2Ud7uHmzwwWkY8uctK0iY1jzwte2WLN2
3oM1u/rWsOqP0pmjMIxwYXETe958ihNi9AX1VnUD8XoLb+tj8OBQSYSlbQflyABK5eQJ2xd1VlMm
MOCf2wvaeBiiPWiN9WmlkuKC/hp0RuMxpCqOYtyY7lkCun8lGrr8uEufAz5yFktfdGvMmqJb/ztN
7gMh/X0qzz8m3kZu61UsEdUV7BeIajjNqRIxoOE7VodYS85tCEGDILUs0oNldqNE86RMgeURsiR/
YWrZskhv9O2IPxdIBIfN6U6o8UDEh0YtCGL5KX7E1bXD2JdrmViXwpjvookV6kCSOWb32u1Iyl/W
LTNX3/GD1JZy4nrL1P4G4oo6yDjM0yB1D4yLq0+tMuGT4VDv8DmV6pw8fzIePyx0Qh4ZRNY8j4AF
MHtafC8CEZhx3qfK8cvp2KOvTGovtCldcWDuyo07j7y/tsT2ng80BMe4FL8X4KrUeVROzXb00Y+t
ddaWD+p2dzZfxI0CSKDkoaKRI+66JgOWK2swgxydcVKhTm0oerM97p57g9wIew5RXUR29ocsMGuW
JSc5CNzSBQt6BtNroUUpYYdEwopB+JqmDZ8cDeNcpSOnPixObtHe24jab1uKq1rXEk6bl0D1Pphd
N2mLvRsNvgRL5BagLfTxz0iXVGqrwtn3e/THjGNo5S1oOBBLlbj/a6N9LpIoCbkwinGGzaZSJT1N
xFJl+f342p8/Itj/sfP/clmQ3qo/zlLSKyokJj2uaGpqKT6Nq45D4jBIpuqa5Dy3sZpBug7NxlAD
lnyIT9BPPC7W0gRFN6g+SfqYybi5l1zvZ2SBcg8wcLdITaSb3pWEl3Vsp/BRkFv8GhpTJWSMHQba
HaDZy6rQuc5emiPiQb7GzjwLfhIy/PGPfJBJor33gv0aZALrAJW+TLkWqXblNaPjrPU3EgqfjPR5
qo0hHUY57aUiv1goyQKXPgcUyhKzKyBL6yuS0IiSMaIAo/pqIg+ilSkGeu5Cm8bJhmQJXPs8u+0O
Z1oIiey+jcc6/Vz9sMdMY/ps2RcxeetBM4RHxkhHme6Vd9daxRXy8s7iZqXH7FNJAXmoQWxClhiq
gVkStyx7O0Q0rTqbgkO/2lt3Gu9k4bSyQARGtvoouo8KuW6Cu6arKfFPaVy0zH+ELeomZ+zDDw8Z
f5T3W/B8ZzSKI/fgb+i6Ip8HrXnnzZrFILIPnFRj4hAIbnLVvApP8knQaQ8pNnEaX2PQCVw7xVm5
qIFqqRMVXfi0ytNBWGZcXG2XsLOGHgjQQyknujI/u1ZGcGPysC4U1DLBihUR4wpa34KOy8jApe90
4RlbNaE3ixwTYYgtd8EAFJa0eg+q159B5AV63Ky3I3JBHZNio7Bjzbw1kq8w7wJ/gxjeYcIlrReW
iVyzAv1VxOOdISnNO996IHiQ455DZ+bP1iyN1yKiYWkzijc12VzulLoGEMUdOBQS8pUhyYvewzTS
DaQpJk4XXAEgcQoIENKcbCRqkWuto9NJiRKqRdMkwfFJ2yqj2vNTU5HPTulb4CyyjS2N+QmyN827
1sLXuq/HG2XtKrv0biPMB5DpP4JgrJ6ZzdAzdO8ibNnWYXspksvRplo/8wFu4rWOQif+0bLdeNWa
B5I97CNMKUBTc6uzrlhb3UAkYnhU4JANNqlOGRR74dxOFA63Dk+N/SY8cxUDFuuhvf5ABssw6qH6
2REy8b9klgeuaF8wjJL3Wr41ZRVYAAv5oPiptkWuFfs/uwET3M1+/3r4xlusSEX2wcLfdT5f/1lT
cJ5ORisAoWDTdnMvjvpyWiwKiveJBz+GZg/kE0NCmUlKNkUCeHoV8KFQ024brN+d1sMpVxB/R518
NH9zV0Dtun9NQTV9TtFYtGPQAdDZfmP/NABLQYROcx2tPR6uUMZuadhsmgNbXwWTbh1Yi0SGUglo
JDliUHZhfDkJkcR8wtxAkNeugmyoVE5zHHnDPzUOeVtihUIND3EsYT/OJOhpF2MUv7lWKLmlX7sj
j6CwvWwjfcK/+L25XvY1dzDIf49+pc1MoYBZzC+Awn9aXoB3OSoEaK2XQLC7uG/27KvmtL1eKQ9J
rCG7yhGD7VcCi7JdOihwVXcQvJzIGs4qxrEWYj/EK+daJRu4u6DGpLbN8ImMGYcH/x9DGxl4/6M9
82mawttKu3kNziYFFVayPDE3qWy0M7kIRMd4a6Ad7II5Ta1QvJjKXb8W1FjjaGUZeUIEImlVHIk+
V6q9CHlrlsyg4HgoJtVWv4OL7cKi8YXV6uqUgGi+veU49DiBoRLI2yfsJXDZFdewHkA1zunANLUm
JR13ItWtxVU7fjVaxcWnd11XUOw80CxoEteGV77wAySv/RvVJd4Ek7/9WiTy+zQQ2e4RBEh3fDCL
cAKEKJvom1RrrDF0fHxrikR9ry6nZPs40poPjkxERlpxGqaFUgs+TKDDRu2L0pR2S+10wq6NHnYo
dzZ061XaaycLRUq0EGZDya7+ORR4EoGngtEyvh/rx5KaOVAqBUFfRkKmBiDHrfJhMCca/33hUN8o
Vwpu94GldYmlYbPgk1PJWpmaywVB1SSpNzJ0Qyo10T9o+l8gaTgrGpWgleBAfIq/p7q6lRni1sdQ
faiK15o15MlMJmmUyuAbYza1/p36bBYvCJadBLFWvMRp1MXiZxNTHgy/P+Vs3+9d2gVKSFvF2OZB
cyie0YV4OLiDh8axJNTBbxtCkLzjYBwk6PcA+Wk9y0owIBG9iUBOAdTxafqdnVMidV2uNqcITBvy
TeazBNczaDULjHdbmYYxkOj/zdqUpGY3VnVJfkrG6XQD0GFPBjcGwWwEYUitfSsdv6L6wF2D0NjU
OwhNrUHHQuv4gEh/6UeVkif7rD65rGqwYtr67Ha34HJhiLyJ/rRGJcXrgOqnvTh97LxXsgJeqS3T
D5HaKNiMTTd006PHi+g2IFkM2UE9d6kCgjFupSAcjcg/NBXBNuDt8G5rdlL7qmz/PYLyuwtdBa1W
Yt8t8PMlzby1apT0tuVgsWtK8b64jxKTVZDYeTw4CAy/r1vz/91HYVsju3cx3e9Q6KV5HYRrgYeA
xnBAnv8QBpb1BnEkQmmsvHpMit9N2VG5/ijmmnjqW+dOHH8M2yPEzIzTyynrNlve8+B6xPiR2TuX
sT7tSGHdvSEYQEuinp50CTL5v2eHA0DQzVKpvq47oZajqGbralsjk37ESIkHfLjIrBqiHN4CXtMC
6KMvLliL/POd0mwBF7EJAk0b/N3R0j2JMbmXOvjJYA/mqwu/EXXzL0gNd0iBTmgYy3wNqfTE0iNV
Tv9TxAv7xtqfEVTA/iEh9gPC37Fbu2hzg8p175Su9kYeENSOZEjwcrcdKToMgSvlubD0GUQw+RCr
Yq/9a0J5s+5Kl9F5SOMwrefpbJK0KRiS9ro9f1t7DPlVlWCDaOypGiIHA98vhNVLUfzIdG1fSi2k
U0Q9pg1q1PRIaxPqAjKRzqBryyJoKBw8fNZ1SXm8eQmLhFOT6tSPPKbgdkOcL/a19Vrd/vw4+nLc
eZSqY7NtOlpo7HI17OOGlyROnh0BqQjAxTnJgc8LBCLJmqLTOl0VyIwcuLOkmmd3f4XhsOCNn+4t
4t85oqsKJgEEfhayoQlrnB1LYNey3H5pC/HU96utc2f0g18eyu2DfJdrH39UmivKbrtg/mMo+A45
SBRkiSaghtnFtWuVgz+kKbfX1Gj0FyPdcjC9TPQy8N7pwYt6MdZFr5fBQxImoxc7vNXhkUonfep/
ndIujjTzNyQT+fuJfNhigEOSUfVwTGgs0J9Bwrcqd4oGSTkT0FvMzoj+BvFk7MO60JEQY5kBfUas
UlHzZ+ob5/2MypMx7Iamn5BKwgifAMJgrAn56TaJRgxvCmT7UD8pWT2AGLRe0Bun0iJODAhNnr+P
tvJX+Ndn0H9ZCAoLNDybi6zVTFh65R/kc7Qbli0KB/3Q7cN2ufu9COWcV567ciIZ3sGnntTggSbO
DDPWhRQx0eCLHFMlgZ2E+P7AOgWCYJpYlFO/oI7hghWp/ksBSd8xJ3hhhh8ZIBgFAeX1nyQ2NF6a
CrlJSnNIdAOYlRWAAcPdZu4TlkB4GzhEVVe9WvfOc7PWn/AoIBcdV9b+q+jKdSfyo21Hg6hWdsGL
s+/ku1nU/pywz2PGfO6dRhGSO3ZVI+wamaF5ntigYXrxKNN9M/FwG+Qq+yl1N2vzFToAPcXv4sc9
6B0MQ3f/gc4JeqzW8+NBMvaoV14/84D72xi7jHe0TmlQymV2fAIz9rQ2hAD4Md1zqKfUrw0jlbpl
ZFhURme1wyfz8D0jBZjgxDQEhyZKp2lP/C/NhzZfHiUk6JUU4IqMqbdmgrDPcVYfVGC9c6aiJEcN
jIkSjm+FIWcf33tpFZ5jA023gocKrd6EW+NgcdKni4Uc+tOZNCi9M8XMYvMvpZx7IKkov+lmGPOg
b6YmL5+ePtvLvkdo72QdSSN71KNcSvlBQ0VpgUbQ9ZTo3/IRRvcgRRhxgQ4Zua4H9ma+1jebVndg
UMh352Ga+guZ/Al6F/W2vYaxFGIPkzXoyJ1ePDzKjr42qCyuSexqnE8H2BH/LHeR9OCSPrEMt2bi
c1wQOZcHuWdPLG2JmFc7lLOjeurVMda7gxH43/WHeWGS5tvn1DQv4utxjkXhtXt1TJW18UewYOTI
7FPnm8K5RjbJOq+Uh+m0bF4RVqHB+vEeZTR6+JkucI6HrESZc94xOMGRPv+wD2tw61qRbxlD9+Ns
X+06kAqoavHEkcgd42uo3X7Jozqij7grllT8neApPwf+9KGuploO1c4jOVVeqZMMlldXSo7+EM5K
NqN+rMMzr8ZA0a9gChGcfXF9YejcSBNfBMaWwkUHoz3xOlZJtTm4zV4WCYrhSayHyIBeAWrQUgrM
t8f+FNOnP/ZdYz/tfQfJI78N5bUhmn1X3a9S6KCjed4jEgaL61lEbxhqNWkvjMO3opWDnHT7tvR8
m3QJBW5N6vDTUfCM52ooEwCHHdnpEhZmZHx79InbdbAP8Ll2K1Uc/6IiVyPY8Kd+xVVnVGACjlvF
WZfFP7jJXiPuNLC6t9K+R3NwpsD9nc21j0/cCV81jWfQVSIvOhs0mCI8/+2kQqC+PDCY5gUJUrRB
RDeNDWNRtCcLzW8KJrHAcT5mn3pw7u3y4erF+h1X/toIdvUTtI6HYsI+qOqQRaJVPxm5knT1sugW
x7bBHP/z8ow7OWL3eN09mKhZoPac/Bgu3idJu10z1lQhKRUtIXAb7PA2FpUuShKSCSBT6pIy5vr3
GDCaGZm+9mhvsLhybGh/X81Wjn/vhdZ4dAF/RoMhGoR05pLBesWNgdt2A2vEfEhWOzfdWCSaxgxz
Ww2HIv4n1K63hn8UJW475o/sTi2KMtP8pPZuoiVp1bmX8qp6STlBr0cNTv8A5XIJbQB4v1+1OFvk
pBdioOYFsM7uSFVwailcJ4KZEhcXP7IAlTVKPBxGuzFQGtehZP7QXJkb9QYcgDaC6rvAwVCR/K3b
XiuAeHEdvCowXKCP5kcsnZRwcFFDGWAvFTh2v0C56goQNn3b24jH5X3DmPFb5RvUjJdLF5vMtJRR
gxO9qtHtAwaas69Uye+Axa4lPnrG50vb+k+Khc2IkvCTS1JwyNQ99+nPS5ZteOrpJTfPlXgsnOcK
WiHKXFFFLB3R46YvBwW8tX9ncXuK2/A0RFTc0kB1m2W3DknrhwVtvEnWtWZnq30785DiZPLbyUDG
y+hzl35iShKQDgfq7mrDSPC0dxrCQ5nnJuQTVGN1087aGMmz02R8gCmUyAKhJ8e1CrF15Bs7ayhD
PZMRdIbe6U9EkXcjgrXg3P1flcfRtCQMuWAk+NllgfWp1dA0+Qyprv6LnDqWnVpfxZZR25CKcplB
LnvdEz9WGQhDJLe3Qeaoy283hPKuYUperwdLWX1M8LBmwSOUE30rPa9pPyi+ye1FZYVmsL3n2Uis
xfKYlPAjqarhRjZfjKfyZAJatykjNFkaomn1pa/maWL/xQAbh6todPBru1V/KCZoFyJEBWeztnZj
fLc4mcXK58CWcRTXcbmqgEbZ/UKQfhK4a87pQ0EFVncYPNXwg+TF2VscXpx8iLv5ZahhyqVKqD7V
8tXOtJzZZwPbBq9FJMQitRJBiqSACyqZ+B1oytaDcbH3RgL6B+o5U/lokzgkccXGY7qCsOj3wOtQ
Rk3rJomYMXMwUeUJSC8POT9jPpI6Aw3yJ5wvVPzYjIptaXpSV5eDI5WqQyDFsvshRc5+gCYgderJ
Nm4N2M2QSkD3zD6txFe8Kxd0DAMdOKJeT1XjVKCSoWzYdl4Qe3NlZ+tBeqLLnUyF8cgEYVwbaZ2K
whBGhW+QJlh1+yivVLOT3FHlo1bZ5njxxZi+VBCVb84Asp/V05gWRPzgitBqDnOXIf/9FDjUdLwR
d1jU1mnMLearqigcUHujvB+ABJy+XLccN21O2x8mPRy1C4+nHIVbk6dXco/NrrAj6ISUtexuXR5f
GFVZlTtcUm7HhKqoKiAFk01FB5z+mrbuS0zeKlrMkd07+WZWzuQr0aRhS7YhYz7rO6Q8iZzvMN0t
oD7Z11hbCacHq7cOLelYy5gkJq5swvc8atmT15GZuWLB/6B3l2BdwUTyER1NDWOj2pSM464N/OpT
AyiiAjibUsApiCb8RmGoH4tse/hqMWkObY3a7xtDxzreS5nXIr3+oQi3q31iE17mtBkq1kGPP6eE
/AHdMdtOMRmQT72l8VID5WIVKWu2WS382HY8FFOwFXEitqFDrsJ/Q43fqgmhvNcCdWYplp4SNegC
eV27HaxpuHSGmP1VYTsxQ1wUS0HOykrQU1HGDmf/hEGnDKsOAY73TQKEi5dKpmHYXP7NairnvmkV
TwQuvkELA2HAMFyjnB+xNsZ2cfSWn531Rg7HrBODjZckHChfd3g56eqcV80msfvmYVrOKFeY668j
UdYbsv2RTnhskTY+x+bMJBVVZHqFa9zhf4mRP6FbfthDvmtKq0rYNgJDqyNQMjm0SobmhmxAd0M4
kIE2LSKau+aYgKOwJPg48KVLJoFjqP+amC/AvfEzpZ4NVgGJdJko/jVzfmNDVEsvaLnCsFUAbUmj
OXABeMx1VEH88bkuqo2jUUm15vqZaIOFfC6y2/b2bz6XkHAmZq8g/dlxVKGYoSyH3BrtepxcgWEx
3eA21GlpEXSxZ319s7d29xPJXYg48KGJDmrefgnar6hQhyueFBq9P4AO47ukaGip2FHjpyqvy+PM
3bNWae4l4j5uCmpOT8FFloMCZAN0+hQY2f6AHY6ctv/RMhJ1UKseNpTgm29GPCQ3rISWlAnu7ua8
xauAN5KrVLnV/a6fzRJcS9estPenw74opiQXuuemKarm+Uu8TIUBYFuXKMl2ZAu9jZmeoiESKnGf
64qWVMiAOFKiwR6biTviVeAKb+gqQCGxl86iqIHOlGVTh8/o14f0VBZtvr1lhzkwjX3t8ZFirfBk
LX8esNMu8+6/0M/CX8A0Nz1dDI36qGF8yteSc+sZX7kGsOVGssXYEFLu79dkGmSjfukMEyrw6quZ
3NieWlvnXNw4av7vBj5l71PqVUMLbK1WkfQ+PB+ksoeeySAuwKSOWJRGTrBJ8OIigGbnRsSSEB2Y
barPjgtEru2wAJ2SdMxGMjb/PuE0XzDanISarzrZBdjp/T3OZT13AI8tefBGSs+22I2nJcNSnfko
4YE5sEsMPq9qO9tQnXhwik43aXB9D6wtAMKH5DOFlf7voygmVMAR9J79TFu9vC8yQkRNrXu3Wa1h
76SI1CyHbtE3KF5dDvyMQPw7PkMCPRP+sjBN4p1lpaWuZ6W6mI2+2zFhRU66eLVFL8EA/OGJyPi6
DwVIZlFiw33C/4LqOtf17PUY0TO9YMZ47HSe5Kt1RotnVe25Q/Mc7gKwK1YY1VF4guoG5ro4OeF6
6gjk73woxLg+hi5WBqaonNaLzczBhiHiFWIBuH90LqEshwSxK0dpD4pkC7ibFNoC7S32W6D+qXtM
V6ISNFvRPVOpb8B4D0qdA/FoAh8ELwIMg/q3/sPV/EfExCtdcZvNa61C5E9a/1tHBSOxVwcFFJQY
32udws/+ov4Pi0mFzWEvOaN2z2iSFM+4aDmShvHeCGiP5iF3O7chKgWaidsXaa3m6Tb0QVrhTkRy
m7heN7WVTROnpyEwrcd+uM5TyXsN43ZzzY5k4Qddf/8PXUU9O2WoOLGmYo5FsRAIr/zUvMiu25S6
tTDeUB87KLB8DJM2HTKZcttKPY1Httn3btjZsN2UCWHaLJy2sEH7vqb0gCJyqxCwame7kPhgJQeO
Ew9mp2/g6qd1YZASGU25dedI7vj/9M8UT5gbGTj+QwdsY7H8WVD124kaBXKexY2htLe6KLqEGxWW
t66g5fF0TS+BdpusYcI3czC0pAWQWKl/e2hKXkTxO4yEhnGjRNJn4FyaTLRB/xtUhBQa5+Tyn8Hf
DPDWEq0DtuIiIYmRGs56HcVSVLk+6yminDL11bFykhQ4moUVfzb4iXO66YPbOism0HsbIOr/cKiI
cJQ7pvUFwbasaE1Fm0DJjywKydqJats+g0Wq4yQDa0i1xMj0TsfQCAymhFjGwslhmEfwMjdiWlEo
AOXb+Kp1hCBkrIUTn0fWxiw+06eop6uI2wdDu+oEM05zkQ9rN9wbhldZAZp8B7zHzJVRmsXgcHEg
GDgOWyx2B27VA9n7B8h4ewmSXsDDqwjx6PS1KwtC5t5jTE4MtoJQ2G7NDN2Up8nCKZLBp2H8H1FG
ZtJXjgDMWQqZpO1+b8qO/ZpsVZV8CmA+2Il0CR9udX0gHxTgdL+P8ChCbohhLpvBJRvGGrBd+HKc
XqoS1/HzIGs5cbWEt/NQ/AsjAAOrMWyG3ghFvbjbPFNjwniNLeyUHPyRFgVqgEISyLokp4o+JYNI
QIFB3kgSR/vZr2Jk87Ehf8Hc68psbnEdq35ne8y7nuSFAvBYIzYSA+bbkPbX5sb2KX+PLDDyDbQ7
swf9KNFNlRwteKGN5m/2kREC0iBVWubSdARg95GSNEhr2Kc61PwGBbmR6UITRcgR262yHWQ4uhRK
AYxOtup0H73wCdxCgXPula4XADkZE/AZQB5zUphXXzu82ubauFcKiwNxypW3UVNcsbzz1kHHWe8x
xWdoPfD7yM7dNtg7jr61cadgB9qdw2PbYKbqDpz0l0SQxupC+eFpJp75xFF8BbeOumRt1ltgvYaO
rQjqxXnomuE3YLQFO+65N+w8Yfl7Cbm71lFyIsId6WZaJFluqOs4ilEISt4Olw1kWRY3cQbD+fbb
U78ALCecLB9LgcsZrYVqwkKjY/72GJkHM5JkWWUSG330/liqRl7PRh4u4YpaIMYuWzNNxodsxUR5
mqdXHR4y86sSFxHb1SHU/XnANUY44XozB8NEULqFq8k75ZBHn/5AlDWM5alhKvtC68BvanJp9ldw
t8MLYhQbNIUlAEWKzL7S/q16evUfjiObLOQFR6KkMpeMNGv4tzryOlPtwSGFR1SsGTClrXXRCOxU
MTNc972JcqjUAn/oKdzDUCD10Ljd5wpT1Sqf4BGo7G5ppKg+o1JUJK80wTCuTl0g7JAqtk8OwRZD
S1XschjUAypbB6P7eaKMpcfOZj4ogg7Oupx6gsgydbHCTI2yRKOIq0WuyIY0vBID4VfX1V7BqCUJ
99B+ulFF8M9LA0oSdLwGaxX9aarBlcvG+s9H92h1/+VM3KCS8xjv7SOg5++3mrQL08kjfbfbbuD+
yN2WgfegFYnLD/+PrDxBUK9xluUNxkNQwGWVgwAIcGwtCmq/JXjuPMSaTSyBRvVrfr7gK2xzs/KU
UOC7HNaEa2pGVqXOX3w2LDJWstuLs6TnDSRgnfJ9pmpFBJyuxEykFKJ5tHyPdbdCK+XNTfSsrWzw
9HJKHger2kknlIwo4L+KFSxALA+ks3yURpxP0iA+n+G46BHqXADHoSZqbEWa0l+pI/V7ecgbmPky
Pef5cxV3z1NkE1eQ2xwJ3HnbILPaDSt0pPm0yz7vLucMvjtD8EmkH1hZoPZt1VBfiBp/pYIbLY7g
Rcx9BqT2bmRajt/cos28PSi7B2hmyX5u1Q+lSoaEPQYYEBZ4CSabwiMfwTpHYT3FtRoHRUBM70zR
S0b2kNhJjTi/eWP1as7r5FD112YkoXWNKOQZ7LlzXEgfG9BEA7UV+T1oCSEQ9AHPdFDdbTjeiWxh
8BtxviYsvoiv9rHpQGnW3cxhS3PAI1GwssNWNlN4IrN/oWdUlpe83h2wNlLQ4ZEaICTazv0tEFTH
JHKLQ0I5itRTV14M1p99hGRfIHon9X/CE54NvhO5tvxrNf4nQA1KRlo93Zk9gDmnCRxgpWuVP/ZD
pm60At+Zw57QoPIWcnn3j7cMqvcl0NpS0aokQuEWtXDYFJtDNjhjZPK94JW6ae+k39O6KrjXtYUn
jTMAmGu7+fq6NJMnpb61+p8qmKEuhrnjFQJ3G2x3zGyZ5yk511k+Ouh6KxFeyodPpWCkzwrSxq3b
gQyGsktrBMjRull0MZgtyyuZVuCfFAYrOIxpsX6RLxMrZKF5aRa3OSpFp63fU69UuBV8QxepUpJP
YnvSN2WS4ymfrqCeMbBKHZXxZctXHBOerZI9abAPrZFU07Dn60gW+XZ7uTg2Ieyj8tb9SvblznAW
vSvxPRood4w64ZALrcEBhdtbuxw0u5dkApRbuIVFOm6AzZhTAXFgvWLO3/w0dRBGFkmkTJD9bMlG
b3IndAu+M93PdVxo3JBL8+vw08Gz0Z1Oe5rp+dLSO8aIuDrlIVhds4gvYjc0GknQ64Zu5CeePYT4
ZGT1aIQdCa1Ra/lDkF22RX00MqpLxt/g0hrtUI94B1Vi4LrKUk8hUMWAzh/5Chfumjx1DCfmFfxN
kl1247IKE9qGjufYFZrUDbLmDYWJXjdJWhTmbbsPM5pXforJoPrWmrZwu/QZgYvI5JrSjzlHxv1c
f/fB9DVwAK/+Tp9g47H0PVQ+13UTDYWqMscJrTqQIkwMmKRjXWk5ziKgezOioVAhZCShZ95dSf4k
oMX4o9/w97k2i7AIcL+1GH97Lz0T8pmUygKX+oZvrQgqInG3dz7kGJNa8JMAUPmZXU+Mms30mbab
dFFg76N17V3dUji1BZgbK9FjEx0dYfnS0lxdcQEHGjeIDBovI+w65cA2y8ZX5IBSR4ZVEo0un0ul
eXmfADnYZOITkQDtWKd5bwkAbPdo5BZ+BpOkFMen/d+JfvxvAgfXBuuS2Gx6wzKm5TtTvakMg/v/
OQP2PR5A9jg66Hhs4gj0FY1lHv+REisHsaUI/ohhg+N/jDjsI6Q/m7nY+edPg6kVCOmEzA+lSHrg
G7QPuWZ3iXUMuyhmmuRBX6GPGqTChofSbIlrU8kledVYUnFW1oZ4x9MwPvzsO34PllDn38DwmmPr
Qji3+hRc+075tgrs/R+XubmxlJv/yVIdIYrNmVXs3PhricjPpocLpBIh7JJx/8g3kDKjJRXSfXM9
uNDKhacOugCUgNPfX+XVfsmJl4lbVvclLpZ8FYPm+GeJm1YcsB0rJiZDAk56DUX3ZOLAvxYX4leK
V62SZM2CtLnokBxUr10UMiFttaf+nCAuyyPLBhlHxoYdFwNtJmpg8hOfxIdhpUX/pLkjbdsSVv+T
LSnwBhG+UsQz6I4S0AG74UTPGySVjUzmlZ5Fxd/BVIWigCB9eh74yrsipXWr2X71oOR6cKJBlpsr
pHwhrsP+ycqhUaUj8heSesQcy2DQc5ET8J5Ib7C/luYlyzSzZFW33ULXkPjKJmKMLnQaQ/rB6e1X
zjuqN4uvwtGdRfhpZ81NvkSCV+Aw6QAR+I6G1iBIsqBeiEzt+UrQ9SzjDZFETBNa0IDV47bbhFc7
2DLaBpc60Iawd1bC/ey4jFXFZvxbKgyfffvKFpJb1n+IL1fdwCsyX4w05VwUAPyHB7tD0FvDMDte
2GfyEM5HVsKeEr6A5ROZbMLVPKQd1VIru3erAQSEpxqLqM8tf6kLTsWkdgY9vjV8q/3b2zy7iaQd
NUmL/ASC6bMVqW6AF09xTliGgmjv0AS9gQanDvYdO3c1vqH6DQHGEabNQl7zSE/Hg3mxMn7O7X6C
FzMFNT+nVWPFrbR0BDNhIWA3x2BwEvMjEkidnxo5xQm0u6wP2pn9aoxJ4MgtN0e5ZK4U3eRBDQR0
AtC5VwbAxxzQZL+pffVubD2q7OF6L4rvDRdHyeWh7d7aGwSZJnD2HQYJ6597+DWyq5Uc2XbTSk1G
tbepS69s+eNXB+Zu5W/Ox4gHTcbvJVv1XiD6qM4nCO3VRLvujWyDNlkpwPg/RcrP6AHzRKmkhtYb
7hO4uTFtFXp4hmi+P+JjuOItLagsApkyWhRfVhJf3C8ZwgKeAK4QYtjn7P3IyEQgliyp/QWv7x4D
Q+CgRLt/1O857HCizXB/gu5I8a8qo1H2wxeHypf3UhzlO1Vubr6UVeryqda+arCtaDalWVnUdB+e
ixRB8JXx59yrzZ5JTqWoV9fGWNZz8UMwTttRYzwyBm/isLH/ix74OkSj0ftttFjh31k2tuOHleeX
loTteGl4TfRQiciHu4R1eYlv6YCAZ74EkcqsyyeEGmXl5tnkv+UGlhBy2ErO/5BEyDqyRe0e0Xlm
Bux0JBE2nosU3k8JIKdkp8hVAAOHvdBnKKKTA8ZniMXLD+YsfH8Xw/TPvfbUES/dDfg7wjf6TzA7
HSlKoIYOZenaqh2hpylLz54WR6YvCqDX+mD62geeEsaau+8+kQNNBttHJtVrYr4+HI8vrNLiAkbe
Yg83pQYWqz7fSknr65hBRyg2pPVUjyWSoNQtkExAdS826/9LDy8jv4Iw8bjqjaWHj8oikkZEYtjF
sC8Az6jYd0zpoycc2NryQ+FO+TliWTpDVrzTl8Npt+gcl7JR0Nz2WEln1KPsmPK3TwtA9DkL2vUC
7upQQXVH0NiJc2tJ6/I05MGHPEC187cIkEWbIG9resqly65YlEuu2L9bhChQlHV7EBJDDs71xLPg
W044YJl6l53eJsbvJWmyDOCKNGCP+jFjylnHFUQUn6FGftJr1JQza0jbNmaVZm3Bhms1V0VeIH+P
QvEd4ViW/0CEOCkUzO5FudueX+Ju28AwcpEqGELdsX8N7Dvng9ZQtYGDF7x3MqgsHc3ZXM8TLweJ
gNNdf+KI0jof7f/2hldRtQK5XSnL5mUayxrMcqfgvY2BF4vljm6fddX1bREVe2zoIpmF3n+j8Wq+
AGDCPd0CBip5jlZA+nCdnUE42TFALm3TGNU4kC9u3HUK1njmiPGj1SgoL67V9/tC/6xtHSu93k+S
VKc7h0o1xdXuQ3YxGxKegFqRbme750FhHLabesnyB1ziWnrNjVOc/Sj7HmSWgqEG8Zyz/njIgOBx
1YLFUms5KQfcbQT17kZNMwj2eo/ObBhehjtowDc/ylzo3TMoXxP5R3qpHm5+riqtfFWNjCHOOuaB
qMIA3ezsHInRb6BtueO/dszdmGmijvSeHuWa75BP2xOTHXg8ZOc/wq8XJ1oOdINqJb+ihbWITBgS
M0k1cMl36J+rglNJ4V1O6f3Yn06e2NR1DeEhgepYWIDK8tS0oFQkozwwU0bU6jiUh7Ao50SMsDIE
oX0OqVRzvqKZxoSpVHiv4RS72L19jXrAaVeMIakE1K4iyHSVs9urO8M8aw2w6+39MbnELzqadY3I
ZmnMQNEvEd9vUOvJvbGBO/zNiuokbOTtoLKdxd3MOf6ywI3Kar1KTcwE1hT7hWAJ19liVqciMrcz
6ckeLlkMb+aqZZaq+Ye2Z2ok1SjBIghsT68meyHVB0eBbWxdZQc0SgqPe0A2eLjwSpoXkginid67
fFMm+b5LLHbDDnuWO6PO5Q1m0uLw/vRm+jh9I548opPLeA4WGSNLLCXWqmlluO3bZqcqVai5JFjC
F0p+M4ePHX2GImh0e0CVaYj20dcitDK4BuKEDupdFp8l5VOI9PlXEinm5WB1lRGtsVu/xvaAnliH
3L690/d5lHRXybEusBZsWlG9qQO7tVKqDVgRmwOCvgE18GjJ93z41kE7f7I3XGcwwTx9AQWk2yB5
IZYOAO2QNkSeZBH0em8PfkpDmO959vA0/Fz60V2BpfFW+n++KMc3ofPkn5W7RV17qLCTL5XsxtoS
ViCoq9BYZCZYrz8bp1cJ9hHhKNRlhDFYJOwRIV7/+3b9u2/jWvqT8M01DCQjjHI5hf4b3dOdjnZs
XpkassmRqTvr1RHN5WK7X4czPg91ZXVeR1rGlroG2lGcAFg/AGQecTjFk2SwDjhhY0cA2dvy+/UD
ktJ0Du1JUxoi3vk0ML0M6n49NCVr/nSAUMROnUpXsVEDPyTVZxQ9qPSkFBHbbhGoT5n+oEMxq5bh
MqTjOKzl5CpS81jhYQUcMxRyELaubvaVdXwogMXoSO4JiqxlIUy7PfAg85sxQBvrn8tbI2SHwXOa
jBb/x9vAm+bf0OUJFqpsf60BjagELe042bP6n4Giq2ZSJw7uVTj4SUu8CcMEPxY6D8zurZVmXR0k
slw2LRIK1EH2R+N/cWsBafDRl24b7ycjePS190rIpIISwvhf9aWGk5m9a9IKNdsnMgNMGxwMUTSO
5xcPgYUIOl44cjG+NJJnVUi5Xs39GU3xMK8XMNAzMuaQeeGQdwX8//1aCiARWbxvlVnNLozuORlo
7yqxVeiuajnozxgtAbeXN8Oadr/lCEt8sW90dAtWtY2fDO+MXVM6BANJJJK2jwtPesedXZXCY1Po
oX0XR9J0/Nzj5EbWzz4JzQ3/jYMjeGYHt/iAg1pKxosoAuOpyj1+jFaqmYUf5RsXSIuB1dIDAWqQ
bP47gQXUMmzLHUpnZWj5ajIVbSBLivpc6cPwvnx+IZM/l+uYofqUnjk894c6Zh29ruciPrXr+vxX
mdQt+g7KqvxtBVkYPQob7b+3OQbdn69Q53qj7YRybqWL96ygDv5d8NwuCmIniwtP7ZEA4Jwgf6em
29gEh6yJwLjhqM2IAgZwkPv4gcCRt3j/gEsSRf8pOM+wEk1jwjo+aP7FWlJw3l+Ms2E8b7IGA1kF
fpTI/z4GGIGDLRaX5kdi8YdLh9gSbIGa4VGBFZowIk03mfcdO6ZYTflKbjcwghAL/rWtvgicEcvG
BKs9R1aWK/o7YEhX0RFdWF4bxWNVBywg9S9ss4VwlIWrFV0HUPM9cMAjKD0WbHnsMmCif/fivyCx
4W99pNRUt78G1NIFXVn6qTOMAoqaiaZEnzqn2ikoDCVFHTeTDaWHfPGNAES1T3ymfSrbAHcsKsu9
E0mXYMFSHjTqQFbPM0ti4JOE0avbizvtQuMGEdE15dZGd2IaO49W1nQHbl99J7pNdHsHrN6VnST4
nTH3c7bikEor6uSjB2S71TKf+UD3B1YxGDSHTil+rocPoKI9FqSogs3YCt+wdZieaR4tCMU2JxDO
rqA+k9u/efe9EFo90cSuGn6ADsbnco/JYJirWAOST1pBXDD2bZRg0Q6CY2CrrNaNN8jt4ib9xgjk
HrjQQGfCl82TqQtD/O0bz0Wzhl6X/bhdgVXjaizU238tAzWuj71S++az3CRdyczRz6RyNJIikjJK
HpQBy0OkvtcOu7YIH8tEqXA7qxifY2E6SDVeiyqzajHnJ16rSm2/57e2daT771K3/r956yds9HbK
5kbak6NhiVJC5b8BRAROVENBwXtbhaQnhg9XNy0lQfhJzXgmj1O9t7WRTWHIfGPNaXFKqWpGdXg6
SH6graQp1tFp3119540/JiMma9i9UADS0dgbf9P5ZF/mLDWqQ6EMoaLNfwuutGpBM0HHYsXir/aV
RUV0GtiJ81JfLQd0BMqBVirEMy5AwB3LPIEkCRT2n8Poh3jQ4sbMbW7AL1KcYa87Ii9vaONKXOTj
9qWngj5S+9OEY23yxk4ZOFhoGAw8g12WAMvwOWSsz3cpfrOHA6qqtNEgjH3BCMa3/1PC12MMlZTj
ISXZmOYOaIoLUrf62jUriYAmbgVWoWlAauWbJ7GC1EFqDPAzBWd3F9htci3z7PIuTCzAuBEf4VCm
LdRCwTs/TxLfkOQVp/T21Nt/w3X1Fi906vUKuCBkiL5tDjLKfAAJgOyIRqCRAp03WYUwaei0a7Vw
vzjv/zvtZ6m7AiCuVcJmAnjbXRY8ZxmtDvJ7SoHzqmGLGUOconIdIRvVsOnE926bOntJxKMH5tdV
cG8r2VUJMxw38YtA3YPezbLVej9xio5jVvUbdT+BvwRhJA84ArDPmMSEXJ0Hg0qvXttUGVo1IwIV
ti3AJUWn2QbmVjHOnr0CgyrxhWmFDPY6H8aGPgM0S1JoScu9Zt7iHDanvpAMBlbQDHKvnQVl0sPQ
EZra0HQueq372C+ZKllxGMrasNb7hnpzob0JNVU6HCF4o1X/J9OX5iDlSYh0uLq8p1NNlP/GgaG0
16oJtGI4UXE0ZWNYgBk3Cf9ynsreq4CJ9TjSKfyW+70IqHrWi5dg0udmODeU7+rjEaqLrBBs3yPP
cNe10925/C6U05okLwtH/+74nDKDorfJdZoto62PnWbrwfIlr+8KXFH4RloHXT4HgEALAjwFL43s
sclSqKTOBygk5bEm3zmxJQ5f2nVnrqdg+g/en1Wb+8dIvPf+mQ3Lm4GiPCGHz48OyklyJo+zkA2U
EiWahrNkjU9dkm0ij3EdgvZN4WZFSKFF9Lyrx39QlrNWc08hycDg7gXEXksm5CM8PjAlxkUFHlGn
Z0NhJ5Sz73DICV4Pd23FpHOp2t374U9oFdzLQBkO2bX0GoCax2QY6JEzb9F5tQfY29HaFqwmXEOY
mECw1+3PpLvAAI4sg7bapLh/tMaTLZfL5BBn+amNk296KUcC+cdAMwQ+X+1x02+In6OEh9+gQyCt
Mr85Smto5Om4NxBrp1lK5zK1SQGr3mQFilhB/NTpvhUP9LzoX8SZoV6Nsc3KFa1t2UkThJVnT/6x
neturjd0JD3ZaDiLz/EEyrUcKYaFZwkQrJc1iIl9wxLkgkPYd4ukiTRR6zzcdaBQt6mEgDMw22mH
F3dn41h9W+5MLdjNEqEhlcgx7Yi8EoiP6p5/SaPGNCwQG1T7CjlYffgmX2/I6YC+NWSCBvaA5YTp
uCNU+IF2t1tLIklAg3tA2AfhcbHl0Mz8Q1KN7RFkeNaGO3v4WknWMrO4dYQdLg15wy4aH4x6Ruyy
PvR7OaEhBYfiHhDCzeIIeEhC26uyVUjBKH17WxnbCuX9ims6FPr1c5RXQZ4MjoE0rLYRtmTnly8x
1jFJLhcOjomFoo1QL9u3tna+2BeOUzf2GDfwhoXdQxn3NRCpYgzFI4P040dmO9N1z4Bd4hGqaSwm
Ro3zWeSybNe6IiftdkeCwXfi++Sx74OHlm2BIS4X4Pdy5xGKoIKh8ThlzPYbSpW34KZIbACJMzID
1S3PsgAQ04Y3TfvvnJ7CHboNmYCJU7pL7sZV1aeYgbBCjFV8FHzxBYzNVTRntg3AonEYTUXbz1JH
Fm/+k5WpD9LwIYNJFdvHR0/Xo56adNcZ0rTOm39kwx3uUp3jJRaQfjPjMsC66pBwRzTPFTn7jEaa
8Rwga2UhbMtCTDEhQfgF/a6YKOUpyq2m0hcG+KDAi4H8R9goEf4VDStkkHE8gdmcZta6LrMpV4AE
mSnrzvLudks9uBHd6OnFP1xLEi670hiSFA4yYr1jSQM/fj7xLuK9z1v3MnqyzpGgUSOUJJw9T2Bk
kvkcwLJOxUl4V3Oz/MLSwoonVv/KptzKM2QX+VLc+TBaq06HCpW+wq+s3VVEz90rEgovplrVVQxl
mAwsLoSECOedlUPd897/rekhUYR6a07NCdG0SPbHg+Mnh6Km9ikMrJRnwm0ZDgYQDzqMFRqvzbxf
UATXQvUNM70E+adCwbkV7U6HZrJdYURckbficgytwWNMxKBEwaUXJL7mxdTiNt1f35bRSkaHVYlp
Gnx5N/kEONfcCgsubBnOkOewubLOymBQmDMzmmBoajd0J2hnO805EasJMyr+LUHRdUEobKDjAENK
kOPgSXvYu0iWfi6Uhc++XBUzK87ZebZlNsNUFL7ejM4BC92UYWAaZehgTmKcMH771Ssz8faHmBhq
bMKivwBy0weONqDpPzfCKgbXaPo0rEs6YohZ1Vs0QyzCeZLoYc2q2vAKTiHzC/NA10kU+DCB11Qh
BAgFJyF7I6K+0wh2NVFIxcyuNFtrfw3sNsnWczaJFmR+u4u9E8o8JHX73Fgylir/CL/ZHQ0pCv+A
PGSzH6uqhQN7pkGRVhwgTpgdP0Bvjh01ZiG5a51WHO8YiSzfOAlkXEZwtGLugi/3RgGUwWvdCqJv
ArJOu+P4GSL3pVBw1ZNO3pR7naYhAZuR/EgTYlPh0DzR4zFUDZuiGCRXvxzaWsOFfFRUJ3En+sNw
pyHSRhn3T5PxbvVmd7fBTDhtERwHy4SKEM79p5N7rlYBoQMGhwUtGLuZrG6ihFynbpYNKDCjJ4U0
aYe0IGyl54p0EO0VRMtZcxN9Gx3aDV0QS/a544BtvYkgu4U5pK2jrRVw4wsBgtVh+zqt2DN9EkJu
tUhI90fM04yUSMqyi3ZgiYraAyPucDS12Wi/x1JQwftjLYZ4vR/QRU+qaoqvH4gApEaDIBuh843X
WDsz/3rzQGzeEEF8UcSRTGS7kWeK0SReTMv/J3WqV7htUYmnLzYB+SAgXb4Ik8AH11GgXG7HVfCE
ZhgX/vmmjizq67OMRrGxf4XW2ugDdGgPIELSCZnrmHcbX2xZJi6/x+kePDZY0m5CNPHWFY03esOM
UgP5wVhk0kGzcQyHzqmBJIqcK6iqP7XRIEiLYxZLnu67AaGH5ObGr1/+0zYPCVrazlEXltsE8cPl
0oljozypWYrgNa493nZ0xwUp0iFflbu59XNGQ4+HVY7xFAJj6qYs4OpEoKE2K7fw0E5SJXHa6eoa
aeGvAXpU3oyO5H9WrPI69TWeUxShA8RB56cH1t0dQ03ii5lRyGXBgKY0sNQGFjDE7D4tCVa8535Q
1wqu4CXd+p1o8Vv8GJw5gWo+8sx8U37Jm+JGBqckLS3BgE1tFT4NMMzkYHOnXTZGJFbNKx1Q9f53
NmK7g7a/x1BLjzfPd8RBQZY7hDg39cvXzaOjzLtK8xxsiDStmacWiyqO75PLZX25PJX3BB7JBl06
6jMul0w5fT1QBDo7FsQHYDazxuDjHW+8mNH+mVMdu1bhtIZJ8Q4fCRO9KBxZxFwK/yvvdhCx5OWI
h1p9VZrKPhxJoU6U4nx1BqlsiZRjSJGTJjLcUBidl5i50k9fFiWLpQZwk1WYMCXp/WlgEQQTUU6n
g39bdU8pHJeZa8EmJr1c+CbuiQy+u5Ze6UGXBOFQT96/Srubyt5Cs6jrSzDbljr1M+nWTeMN+0MF
Lx8d0aJ5BHQcvDJ4wx7w9xBGV1dVVkSdXu0kAqR1Q+WI5mH13PPI+KcwZ1vbp7dhvHUgoaJg6GJC
HqY5gN38oaTHmBwiTUA39lPFjqpsdnX1p8fhCDwAMAATD6IV62ULSowJjO69mzBdTTwYgn2iKJqq
vrDTAySXk8yQbZq1Coj5WB8+mnf+ZUBxRVLJSu8mZjTIWWRaayJUmM7RDOxid3UMbuQ3MHnbjSE3
CYPhkae7Ie9pCJSC5yyXorR+08agJz1Lr82Ih4HumBebihl5lqzBjAhRHewFY18iNhjn7AxmB1UN
hyOGrN/rr33CFah2s4lBQ97jdvesEtx3QGfU67YiUI4shlustQr0jFDWU38jumMOsF2CP1IhBWgf
jYk8Sd4zrYNTL4w95eUJ3ylGIkitvPNQpcOlQgKkXARWhXQqM7JnS7CydhoVsapFzqYp7y4WIQKb
pJOOh26NhFHSiUVUaDYdXrWRO0ICU0ES8wrJn0JW6DggTugeZPfhy0GDqG5GHeMhmtuOMC85sE9X
tQidU0F/IuphzaMOOyyRoWZuiSKr84TwL+VSMH5lfQcRYpc404egIKx8JG65L50Q9C/darQioHT8
SfaEb3eyN536//erHpJTX/b6h5BvyrL9FWBFUFA84zXMY7YjfROec8yj9wKfIw4Gm5pGotIh+7Cm
Rq1ujf99JAnWh33DmU0XmvQPpabFQ+RxoqL//qY45EI4OtiNj4upTuLIVOHbJSbwlL4hNqb2CrIK
i+MT64CDPin2Z70iVNfdKt42q7BwRH4+J2iAEOlMAbbL4GmtyuVEaHjsincUTO2ZKlnl1yw7Wy1Y
yrEULMxj1fBC29+diKF0PrDVi93nJhrHRGVUH1/fhKNdhVh6YqTXbMS2Pu4MY1rbt0UzIfUG1I4V
ces/uI1yxBD8BH1aBsMf/syF0poib88zqdi6+JlBTwvNd/6RrjsjDWYOh3ekMYXsDw0Jq7DHkb9b
MamW68DZsuB9dw5X9uIVLRROeMlTLNQlIiSmosogKiQYBOdaAvfaoBmhN5gJQZ9NdKYjNirGY3VR
QA3oke6BvSLnWIsSXpAb7MPftdSf1MSvsdXLBsCULu8BQCP8MUtpJzrko/1oFzTkflyLYHoQo0VE
1JMZxYE4IAzenOm5xbSG/GjB0KdfyqEjHIeESZJc8T8pOYLRsdLOu2Yy8fmI7GNqO4ZJl4N62EVN
prLMN20kHcmVZ2Jx4ygPnJ8IX+k800G8DuUctSncFQILY7fm89xCl0QX/umBb2p5AM0HwUli1Rc8
wvgM6xqiaC/mD8Chsk0ksIxwu6WOUhyJ+Zn04rMAk8pfGq803Nb/mLTfKaXOOszVY0gLib+qHHZ3
D31IuExfIqRacFGc3ag8GAWYwtNZ7b6y4wtHQlmMejAAsGCCuUOkOsEagOHTND/SQ+AgaZIF4xSy
mpJM2i7W4qN7STnwUKpXGmgiufQR+/zFvIK+8t/4cMo0dzonWBhpMWdgajUNzVa08WQqQhslqngu
Lr5Agj+wCiqOnjzaGYHes6gFuJjzlpIV4xA23W7wsrd6ZN5wDkfk+J4lQlgZ1FKk29KEhN7GgN3A
nLsheGHWVJQ5f4cZUc0iWy7IM96DBcPITRJebhy2V6LhzrWN+m+3ruI3D+glOmEXirNnVaX7Z2iJ
EwpbrVhCOhmR1j8OKGXFZ7O1kifEON66I1dPONFEib1Yo5tNi/XAXqqerkn+UsGTU4D3Asmm03+5
soMaLujsCO5IxXhWs0AoEScd1jhiIp/9FL7ppfMHM/eXlwXYfa1zYWBUDpxjtnvE+hhFSYlC3WvU
ECYAQ36gQgfjnu9taaIAfXkkoHS4Iln0+kfYUVkLJKZ8f10wnD+gBt8ivMMdDGWPkLixwxr4o4Cc
I3Z6XKv8DfygZgqd+Ty90pHAo2vBitk1YebYsKHXCAGnXA11uJ2bJ81+ym6z/YC865y+Ujxy65fu
QJNdABHhT4XcBkgBrqbbvmGcsUD0SNk8e1o+jSoLt8a9s6ST1mmITRSkzF3S80Tz9WeNWLRGZsdi
YftrW5ieQLxEIsO/sDpglQctOhSlWhX4WynkqOX3WA+Upw0o9PuGwmXU5cQj872ze3eLvtzW6Xhg
hakvngVxVWz/q3V27qwEvKdNVR79+eq4sAUNF6JSSNNHioIZLZ66AXFdJFkxw+05Pn7rX9wb5cRL
BCgLEZyzgVNkLR7AwfsEzHwoEuH2BDIOMcfqmy/6Hi/ANkcNAS7d5gInv14Hef5AwCCNKmjgTDFa
wFHJ/lLmu/iAAxzIGkyvzZXydHXWRV2wMQPkcZu5v9hCLbxSoWa+oJ2AGptOLhbxZkihW0pidLBB
+soU7igHCbevbtZg0khX6T1NK2ZKEYk8O/CoD6kYqmyZjgPMFyyQhmUue5nfu46G7PDwTLk4VeHO
s5ieBHXEhGX1KTdpiZXN72h8xAMnUVh7/fD4d6GKyJNrfjGmbawMIda1qsM8XHD2SCwO4ltShRZc
CMqGIpn50KniTBFJWcSNKNbRYfJT8eD60bX1ah2OgBblfSGi4K4+Ec0T5N+ExXK0NNQTRMlYI7d7
loqq6xTH6AuHl6EDME9mQhgc76kN72u1nEB778gB97bevA7V8JcloWUtmZRJuDgp0dV63JHOGwbO
LQACKx1glKJQDG6P7KxnSwfQHMP2EJFQgaEByK6SZnwjYpKUyqy5nYAIPVhpGp6yKNGf0v43i//f
LXRF8VtnI1ng2Jv9hBlKspVdbEZyedMoXv/3c2qahfvscSVa6ieiBT8LSAGLHS3pmU9qV5zJb0JM
73CQqrSmaIeKV1po5dT21T5L8lPvELaqL/lYM2KqZigb+fG1eNsQpzBe6pfItYNBt5c5lkag61HU
ICspll/22CeddEBsfuNJImlyYwwVU+ebQiFUuOdnnSPQix8GyTmG5Pa5MY8FD+ZdrtD/RmGtMmFk
nXWhXUt40RxLyM7NC6ncRnAqtiQOgpuCFXDnOjPiEHYLrOPF2arR6jA3De23mnp7sdaWmqUGEdqF
bte+M5O2L0kSQLRA7S9AAiz9hGx7MU+E6AfqYD+C4kC3qRbJWNAucGrI0tqfkbeZYiogUzeiwsQ+
yT7xHFPl+VfwYDFFe/MsZt0VkCH9fDFzWKfUNy+z1x7FPuO01KLYBblJYfbjxe9m3STGYIXIGamZ
+F8pdMZx+Gs71Cn2NyfRMjhsYsb1AwOYAXlJB+OmT46vp/+keCE0ucjU8zKYD0cCqs/zb8TLqDtA
IxIz4bfWAAcebYV0jlUiLNHIhzWA2UXudSKAIe6mnILha0+ubh4/MQBGlf2/BkCzCEt8hRCJUe7P
wzJP/kH8diSlbfcSy/nSzn8VL+uTa9ySQVnBJCzV3KrUK0IOCwfdFayiANM1OJ6UvY30PHF/V+1o
gkOQv6D8JZ13SfLYWjv9DFfoeCowrgDffktZnxpgWXkjBp+mBU3/GShh8sehky4rcNn3l0MFhkKR
y3kxX1OGM7X1cO0Y1brBERgZWOj7qjLOLewdjVFPa0lzWcXWpDO8yCaqI6PxdNQ38/wOHAefOZcd
5uzp/QP+bicWdm8Y7avJ256Zth9Hmt6GPH+3sVxcbsJ5C1On2xQ7i3V1qe4FLjpF+Gk98iDg07PA
qMfM7z/oMnNp9Rek19KVyEQY+L343mzNENeYRuUE2EdI7NlmlcouyBKTg/F281KPHANPM3294gL5
riznsXXyCcbEiRik39xq0JjJzl0JN6+Dv76X2luN9p3O7/1pxnIwMIWToujbhktRGoVt/0EA6VX6
ri8frXgbQ+eJ3cW+2EetjoCxbHO8d/pmI+ZDZQ/CeC+4HY8MybXj6Q+ASOpqel8USs7/qrOLf5Wt
tlHyJgwASWtPRtb8FR4G+Evo4ErGx96r8M0n8McxJJorSGAbs25FOm9ZKqcmFGS8+3BbRZq5/Vc1
0yXJWQnz4ZuBrmoYtBpOPOi6keJPQR1ud+/LzOIyJ3w68DvlrxI7HGi/KPb2tJ811RtttDJkhu2i
s4d3XBp/piVv5Xtpqpd/Xn3TD0abkar3cBjDCz/S/ddE0F97a2Bql/YidNmAm9kIwLeiGIvofoXB
FPOTS4CHzpmwJLXJUUXotl/CtH6KFD30BRCPf6jOkke0DE8ryHwXJdAT8GcqBnVCwSzF696gK2ea
x/ZNU0XQdQGpjrOENtf2XJxOaxsBp4NUh68xF9/Y0GQBVe5y40YOQ/wVuhBuEA5SuLb9I079paWE
P72wmb07Idx1k/dXAav2WVxBh4/LKxJe9XXC3B7Cpj06wl4jiWfH3n4awRAS+RWcqEJ6FSX9hXpM
wzmPKZ3usKPMi9KZqtCXHaeDuaZO+dipGqCCnq9BH44Ju3n2gVsQPRaKdEpnczQsIXCRIBCvbP5c
BsUDrqGyTZNzA/ajyJR+dp+amZRBOEDRkByAw0M7SySJWk+j+t7ICwc6tKKSKxcMdRqwtOtH5hmB
g6ltO/7niK5Y0MfVFLeOVtP+zAcM41K+VbpPATOWWK8K4gluN+IX5Zuv1lmIO9fKBB7zvtPrtLve
ohFuQvHQF+ZXI65KTNV9ZipRYpNUEyk8WPSe9ka9sxl01wuZ/vQzk58HnHZ0LgLu7dHddurSyr8Y
enQxuMICM9r2hcB3LuT/AjUhfhcMnlvPxdqyjeiTXqyb92Cwp1ysSCpsQemSUVo/sIu3xabxq0U0
gWzB11604lNs/SU85sB3rqcvc5TRxXrUdulr0zbrmLTYrtHp0XU0DEqliZY/5TJZSRoE0PAvGTXo
stLINGxG4Za6OgS1URYEsnaw0kT5APnmzHzu2NpR/w+bj7suU3ZUUbw/Hn/uPYO9MFRJ0DJ2XYr5
JmERoCqmtXfiIPts/xNX48PZNXAZs/ftq+nvlRE4fGnunapoqJ+DyW3hCJtaY2A39MTQLImiyKvO
bYCa1X9frOT6C30n/8aG2zGswqf+cfw/ZL73c+HeaGrMumh4IC0+S0oxBUnVwX+gaRl09N465TEb
dWXcR6U5nfz/7Yp2a9L0g/tKtc6AN8XCqQK8bUOTVnKzar2E1bdHueM6Y5JMjka7yHac8eFL/mUo
KFMDriBECyonH9E+ct/SKR/g8957z/z9VKZn/2SDi5OnjPnsyIM1zTSHaN6mjpO8ailqYQd2nnN7
XwMlSFRKzuEKWHizn/RrAPJvvuU2ri9jzm/R1oV2Ci+YL9dycP8iGXLEluzo9mnu1gjYdbqqKsbp
eBYTrECjRXkM2OVXQEJ3cj8+ik6xadmDHSXRE/Uf7rzSH4FmDkb/rZjn/fn2q8vK3f25kokdTYTS
jSBt5rJNMJ/YqJkFGzk8U3AHzLVUkYujV7jzmWLaSn5Wlwvzs+kxmJusMoUBkwyppjpyaVr1XKpH
yvN03/uujSr/n96ju3WyyO8Ifw5ZLTEHy4a2wmysBloAg0AoEEfJzKbNTJsTqmaXBCxl+mzZV66n
yWbMtym0Pp4e/3c98+4aFBz6VW1tEfmiUEgRK/xQHe3aieZBhKjavhCN7LtZyC/gLgHAeEfPaD3v
KIHMBTcqElbOe310SjdVDG/45MLX5HpqrUAwR6nVxvFY9DyF1XwSbuUpQ3dmRrYa97lX9O1REZ6N
WiGsSKKsEht/X6ydDeAqnF7zp5Ln29wwaPW+2SM+2sLQka5tHBHYHLnOrqRbgGdyuewKSS6I/k5p
+9r1j3NmOoGe7WyXI9Bfr3sZxKMyiouoBjI1AdqoKOLq8xQoznPeoaNwaI2LD0AsNiWDbIQiSoQH
4rTd8L9mnc+cFUi+1EaRYq9/4iwdNTaELcpuuUWCTZeMIQE467e5Fyf8ni/A7lE42rHOJjALypbp
/4+9i1ecDP7LPWjNSQyfiwp6nkwXHbFKvdQsZ/0LnEtoRi4pd8vHt2w5r5cVTaFMU7IGe+g+l7B6
ltbYNyVR5EYDcQICidcabXUECfjRwhnRPlsSUtqXv7PIAOueBY1G8l4TQZAJyk/MSRlJ//rhTYHs
9NRFSnQKCetGG/tnjEJ17Jr04mvNQtMiTF268xNAcyhB40vo/lEWhM8PpZc0hvy56uweG1PZ+1lz
URqi9g1v+Pt2/Xzc8Yc+dbQjqFPpXIy2AAt2PDO5Btg9R01nlkQZsdGyTWp9cNhGaGSUmMhqFwQ0
NbNRwz7hCh86Tx6tH19Gw5oQRURbbYCFcmT61Xs68fznre5rwivGves7VtDa+jaCLmyRBMeF/v2y
ERNbOE/70Ed677gCDqRleSkQKiX4Tgz66aVWzXB+8DgWeBdYW4PH6O4jF6Zu7Fw59UR6EYnUgvdh
Z/6tixoZoO0jGOEC3rvqkNOh0UmAXxCfXQVaIsKEWSs+tD6fNQTbku9D2Z3V2MG2XJIfps7jGTbP
V/RnZnwC+FTE52EEb9u+BSQFgh5hsARjso9C+L/e+PztrOgo+sRwrq6H+1LBt3Q5+8VvRKO+5sZ6
KtUD/jfffdGrBeDi6uAMQgWaUSgLt5V34QsTjT7V/ctVRCu09KZ+tVYdASirZAqkpl9Mv3Lv2VVo
XxLE8GXl0Mic2UOeAMYAM5Y9AY23FnjFDGPXZSN7DyzdY0BYwTB/kDPDkP1dsvqmmu60IBTmLSd2
r3D9TEcStZH+klotmNDbECjaawJvavntQ5uR9iYS2mYUAucSGKRYYd6x6dsa5u2mQJkYqSv0/iZJ
t72jkAqTN0heNTAoDEPZYFTYDqgbPQthVaXiImpCmFuA0GTp0ZZPmp2Lr44DhL8xc7YCthd31JyL
peEtr+O5luLaxcOVssVxc0mhw9uhgeYeYav8zhA7XMOQnMpPIft4YU/m62D6xo896Ka5JkEITjPy
VTvF/VBreO0TQdb3lqzr9rLGlWTbu/CEK/EB3LFn14AbWSu9Y7yfch8X1NXHrLrfAI2t+n7X4663
5dyopMuecTza9bD13jVt0O9n68HS/ldbL+pyCiCM3HZ2MO9d05bCHxwy7i7IE4GDKuQ2IuCS8dvk
P2/oX6DqIYaGEjF5CtBJwhuiBeV6iKt9wAsO/SeEtll9/ClCxnaSsgrmqSEPm/Gafb+CTSwTOrJj
kPeU7AFvjarSafyUV6lZp8doOE8VZUBbvl6JkcjuG90QknjGlM72ANBqYHOaapxZVS3dXRP8LhJG
flFPzRbY/wKS61UWOesYa3PKRQ65hzca14zVLKqRfe7pSfEPBo5J4raz9getME5JoF7RRHws/cYw
0sqV9A8bcpRBIF8lnIbpqMUCIuZD16XOuKanMRBS5l4TVEYyzKxJIMGBfuAzYVnAIn3aANJydMIQ
pUWDtZuSMeGTjHpUZREMlLVrlXw3dNlDMmhBmcuQ8Fi5IJGZD/4IJliaVyf6fokEa6VUvKDnWQ1k
HzUathB3nvC32rFYQTzjnrKDOaDuLyHv/m1MJG6y2RhTUnsJMZZDGXbZrCq+GdCVRmyyP9rEMdCU
rU/QzeYGrMPIV8PA6rFSjpamRtJrEUP2xI2qlw4h7gee6jyDxWsJGMx/pYkwmrdh2up4+IKCQWtB
cz7/rIBNz7fNoARRGEqb2cBAbX5jfVDfjurBVPl5nCUjGKHVs6+be9Glvnc24HOw1DkDCU5aKzDA
C9IHqywEZuGSYDH7wzUgwtqIC4XygcNkk1DXJ4dS9z5VBEvIsjUjgzAH6QAKTVpxvKwwNL6k5eM9
qCQyF9vG3srw+XSGolmDH/A4OJOVLuunA0qGVPZxcKUZiN7ri/NtR42HBZZogiHO4cppWWNLC4Uc
Tt5kfLSYST8/gUSo9zMiai1teATjrMt2Y8TDf5Ujyjd+rPTZJmwpAPuf4ykJk23QWNRKVNhQC7R8
/Hjb1GtoRmZ8iQjKIKT/35P6l4bN2tsaw9gNYIcGhGCHMyCIarnE/edMW64scgKCd0k/IxPMJyHg
qivUCH/vQKxzjgOc22BwUkEN0ez69uzdBgeBy+ht5tE7DDsWXcYyvaMEO/kFr7IbWETuj6nrnDKg
mWhQpLePypIzAEYHUCFNZKpMBUkBzDbf2rasoRpXWalryaRuvc9Syc7Oui9P7bN4zsvNrmPjqwP7
sRiVj4eqHA0i3ln6BrO2aH4dKfAXfTsNPkGn4kudsmTH6qKuHPDLeOjzNVeuQ2z7IvJu9/JYJ78D
eMRzcozSVJEHikfZgKdJudNdep/P0JE9F12SNX9Iw6U4cnsIGHvPJYHahPWIPwgNyYCTbnQaHPjs
XbiHaSSt479YO6MHxaPSJKkp3RqNPiO9S5bdEgF00RVO3ykgvA2qRGUSjxAIGkHBkFKK3iWhHr9T
roEk8+QgrMisE4SYb6vkpFFcVhpQPoiwUEaUxl/awB2ax+F2QjrkaZ9RTSnnp+s3Ppk4cplsEepB
Axn4YNnPboQrTwCeZfjs8/t+ojdQv9S8ZNfDn9h7H1jUAZ4gbdt9qw9goenXfESm4BAcLb94+63D
DPW9uRZO/N2U4CPHTxf2ECH08c1W1ldxijuHSIAK1eTx+oQojv89NEYXse81UOiZA6i689WxPsSP
NL3cO1Jc/D6TZbVfi+WTzLTHm0b1hXWQBcUsfGo/SKT3UDBWI9krx8IcK40rD3vHH7vKgg1SuMBO
41GxOlPnopBwZN1heXDjjUWEfZPoc/1BEihhpIO/J+OcHQaH6jiiDvb0XMjzE96Z/U6nkpEu7FVH
OtAcDeKBsjA/K13p4WEPjvixMQQtwCEeR0FexxfmESQqTzZjDDbLREMA4nVhlHruA0Af0k5/a6nq
gAJpAr9KvvhUz33WVXYqQPU9nocSsmMIG73yDegL1oWwUcP5YjWQCUCF1EodpL6QgNrinz1jNMlF
up/+YSYXTTEEFPQGJpv66MwKzlYlI0Aniovxwi3CEglM4AAlE5h2pYxeEeGHsbI9/W8jIg3ytDMl
v1IyPUjwZaqysHTTnuryI3b78jzdMfRHrWmx3d1J0k54zt/JyEOs5foPWv8KsKBE17owtSIYjAlK
2+3QSE5iLeAq1t72NBACKvYKawJm38LYhyO/1dqK5TdhOkJM6x1v3zpgEfL/WKdqyrZpgwMHXoGb
6wqa4mKvNmoWeyCmdXfDzJe/rM66Ahkc0xxsD0QP+prZAkhkCJlpI98faDwdU8ClOPgOuJk9AiLp
/gZTDg173cwf7YaAdJjOdiQdRN05/bbygnNuvrzjQWgMga4Kl1HAWEA7Lu7pzAS+lSXAlvQ0Rrkj
cPlLV3sNTZKHJVPJ9dangPNJTBMXWzBCTJDNSeRHobm+KjHKLHMYMuhnMhdpVtyPgbNGHBrvpQFm
zf0E4m4YBYwiEnfqm7vAyAlg5RbsCCWzRZuk9yAXnqTd1c7pyP+2rUrLERP+9HrAztiAcPHFfBDQ
hR/ICoG9dUkNfcorNa0Cpgqu+vynaWB4YIPpXSvsEuC9s3FWVanaopD+ceJOVmVNyAi6b7nI/+OB
eDHUweuHzCrXUOZ94K4MHFOkNg6ZiD6Qv5LcBDNc68JQbBVlpzwLxLG72o0AXA+L5IJKXFPIJecT
nxy/AsBW8nyhxpOUeUny9Au4f0AJlM+krkwzsHUq6OLjgyaoAi/4ue6txHYnC5cjNMRYSCVEhyD0
/9aAK0b29opBvNALvvnWoBuatbx/Q33RX7QUXYMesKCu4WNa+G4XOpF0FizIurnLMS2JBm+gwNVp
rg5W4DF2FyUTXE5nO9Ph4dZ5f2JRutywet8AfAs1+dK0YXXhwE7M7BzTKdXLTTrZS7ugMUnappR9
NfniaXzENTyIO1SWkekgfnnDpzbN4xuMu9+fM/40Z/KdzjAnOtM3WOeDL1bKwCzfFea9GR4cf1kA
rjajIWq4tYOI+OWftMObpU8QcTvrKsnlsO6qsKNqNyKhQeaia250+VpKcuFJ1QvGlD+CKCR7X4J2
0UJJqc0o0iCbj7GrZQPlpfmeuNzgBvCs54RgEFbc2QhQ+XV9pOqKuk0dtn+tv2We/TpsRsQHBk5B
04T2tqgYZRFHhTKkYjx6P/x6VeC+hXLsm4aqVQMa0NGhX9zY3GhPT3Dmv4ZljyCJzAD+lS07N87q
cakE+a01vqhLZVurZHyS3MDlvPbUK6s22ykBrFfvrmA2hqPSi1ib1Ypna7rphJlAhR81TUeKbFu6
5+NOSMwyJmExZ+HeIV1CG0YXEE2+PIG6lu7VNniwahnU569y8Dmwux4I9rsACevEkvJTOOOUX8sh
C763uU56ImHCAYxugQS99bE9fD2PjZuD9T0W+DVrtfNx2J/xezbI0bjXDd0ZB9NEhoISBvBpdbzR
nsHVFvHnPnUdMEatJmqfHk8ABR+FDHiN/sSqqBc2ZSfCf95ax68QhMX1G+GWWXBUibgufYFTwEQi
Ro1Pa5Q0lRJeGPJM2BsQq0AuLbt7PuEGFKyTcMW4KgfnVGO6JWlW0nfjmn2V2fq1deMZ7iohCD4O
tKisOnMt88Xw2+ONQU0zILE9qDB5Ax0ftVY297D4oEvf5E9Kk9wthsjssHCsPm1jjXSB6ngRmWeU
nVwp1mq/chlP7rYACeEUIZUqayEfrE0rmnmw69vv1muep2HajNDq52CyaTSNfQG5UsrIqTQhK94F
xwqLWFZv7gv2oCElIEHmzuZxZvCGNYDRDy1366xtalTesbGwNWS5IXgtsnaVF/7cW5nfO2wySken
G/rbjZCBOUXZEIwTCBuzYm4+24drZhVLf9O+gTGz4kKDilCR8h9UxbQApyHqe7ehne01+m1b/HRF
BpGTxCb9ASDzhnYPtZ98o97lJtVyD2TUNGxtuNE9Dmxn25uisBwBE1PBs/DsbRW/+0vbymOa5KjL
nsWRK/IWWewek03HgZ8ZWq0K5BdTH2cqeYwh2bjXE5KxGLejWJpS2MATqlTbSQ7EqzaPbUyWNwS2
8pBHofrM/oB/TvAbvny590fYBXbqUw1EIS0CTi+v/G4KEJdpNerpRPabISSmS7BMizwgZdMXMuXT
DQIuVF6QACe66Dd/PBKp8JfLDbJpyxwrC8lMYZQw4XEgjWjTMUfAIurG62WtbFznAZlGFUhOXDoz
eJEd7ecA+232GeMZJ9WdrxCwoQVkkssVyLwGO1X1X/YVuRGI5nFBE7jsBNdZpIJ++F8Hsx3eUn4Z
4fYHoXb3kbdyKK5jbsrrj74PFth/nB2uJrIJdaMXsonMG0CetzGlegJUMTmf7rAxw3eaasWG5L7G
BVvWdTJYM3uRX9OW5NsyEKe1miUTTRIinTIdFJkT4sgr5a2EXjK2R3PDjIAgEXAiIjJAidY98ZEy
rA5I/iRcr5JAe3z5weOHr4l+nwCbqTD9r0AXpOBeS0J0re3K+gdftec0xguumwQm/+rEmpsMFEWA
oKqPkN3Q5WZPzQbiu2md9KzLCILScQp6mK2IKCFDvim7munyjBLc14Pn9zyQkBhdYXo6JEDdD8nn
aXDptzh3pGRzyzM/RqkENJ7i+KJ7AIYDCgIExHGuLP03FC89AasVllHSdLoPfX3xjB6Ii+ht/qYo
LClCIsz90Te/afRUhP6gZxPPVHzzRyUg2mfv74gh8FD6XGqysyzg6NwOpc0acRuhd7V/yBSAJj2p
s0KuxemZaxYPbwoJd19GYZrZWNiVl/Y7Dy6q+jaZpswp2rG2vv6wGp6QrKuxhQ2yQiGTS/coLa+q
hfx4Qv289P0NK++GYZy5O4z3Q9svVYU+8vKEzGzD7iiswy8Lhmm7o3IsOju+LuudafYkLyrB3RZF
fZeWO6MeUwwtVIxlW3AGj5QHE5cCra0uGxihLgPOjvYBdVx/C2BDr5jlr5PrUsxdqzbucqsH7EQB
yjI1ePplScDv3O9k71zf+SnXvIbZCwLEFce/Y8iHIGTrvTf7dxsVojbLlizqKIsCfQVTy9yFpHQj
XttGnpyfQk+I8+C5ch2GXoiC8fClby4KbyRvOMu2c3ulDOwp5B20rGWlUnI4R+Ws3gTj8VRumEZ8
pzsuXr0qeP1UvGD5qRLO0S5eri0Eynp1/7roekVC2qwVJSswsZBEDg2zqoQBDLNrhg80G/4Jryy+
zqMwWBFQQzGtMdTTjD5rLbYCudhcdmRPtCo59DY0H4jPjhYAZK3wsVJ5vlqR1OBOc5OkpMajP3fv
YidrOZJvijOZtc5LIH7KilOB4hzxIvfGWkNGbnW3Akvz3QA3hsQRRFcTfSbbqlJr0/L1y+N/eeHr
TAVLqg1SRY0YMzz0mum2glMnAQiM4IhIAHeSIY+SlU+m97utzMVcSAj3Ob014nWzL4fat2I2GBVD
ugLlwEsCqcFQMGpTgyylU5RBPy4DlpXI9h79lFKe6eNqhkLoDqbmGe2X2fP6CSs7Deg0D9gELFga
LTx8uExkMvFLZ1kLSHOVHAZqhEacbpT04zci+RgHUq+nFvbmmN/h1SxvPeO5HsilH8zE066vtwiH
nNa9zQKZzZrlc+8So2bOJqJI9mzNq3wukdgRlbi3SaZu+JYy/GI0Z+P5rW6vB+e2SaLgU90sF8Wg
4UQQ/WstjWobjWlWoDwq6wXSixNxrdMSnFoSS1RkF8ismYkXyhr/kzZgyHekMva2w/O/AAbD3X5O
GsBfDoYVdBT+ahaB695jz+D76YX0VFEebp7XtGhiwzR83HI7FKPS+dqkFdqMvOM30lfrj780j6ki
rCJQZYOtPb/p5ATUDlZ+HR/NEuYwwQ0MnVxiYfSEB02tWK8kBR/i4QX4ut75h0lamD6I33cFheGF
AXtzTi5felydJLWe6vGT0U+QIEB+AGu38MvnfFRdmleUxsuPjw0ctO/CB4dVvdQyvvLzUgByo2Ek
03g7LkMBkNn/Bd4mgK+X4kvKmxNteBc/tYK+bRe87yoemRIbe2LpAacFmAUaFY4fnVAPhqI33Bdp
4xadGXvIuo1m9R9p+ji/uICwCbJk+1vzpsBitqV8nr3ZuL/wNOU1CBX5c+Y+uF7vtcxdj5Wec6E7
Fzrg2PqZJcpzTKTJcU/7YOjoRtNYPqljyECzWBTcPUmy5Ryzb1C8rQQiy/ynOQfBQuxv+yYt84so
n3BpvqxBQ8zcjsKpMGbqKpInwuIqQRsBk6NeRVSno/YAYsNTANhKtId3cJlUzBzAxkq37I0OxEZm
H6NaP0qqs0ZTv1MtW9AiQ/7nPHBdRXhHWiBsXxFUBvoHh9WRcVunbdO8ZTKTJ1MVDMl6UzZJ1c6L
vG/SR52ZHyeYKIpFdAMl4tj5RsLsOwkbNkdehPfsRwnHYChNhIxZQcbODF1S9FMsG7h15dNHAhfy
2KGeF95IPrkqD9rbOTdOvf5bFAO7bUz92Q8Jqg1T3C3cK6mr618jmP4kNwCFr0ZwxIyRuAeeNgTu
eGNfvJQYgWTN1FJxsjqC28U7/TJCqRohxzOltrB6b92PiIbozutuTqNBYqOqEmnM57OgqtcG6jLd
0VTJalDBhyAB14J14x1ezPCP0MqWi4AIB8Ew4ueh7+Mh+Rs86QFjEtlvQlmmky6d2MYS0qit6d+K
mh2iI9OKeRFW3vsMMq5Z9ZFdslzsapar2hEqX0ApM5sMq41zbPfohQdIFqnZyj36t6oIO4Wd7De9
cUdlP8LTd6XH8gUfilk+7yks8ERbtPGDbQIc834GOrw1tnN/LKJOmWQfcYHSZWOL7CEshEOb/Av2
q8X6u5nDFB2DQ0yiNrU0veKUJIW99lFk5CZRdNny/OFDgA3kySCLNDmgcolYgO8AJdEHyPyWjKuT
bF8XCaYhWFTgEzsH5OaYhuz9BiQZV+z9wRSOCbODEFx/p2wNWKHjGelPcNfiewtM/aexNrWxTux9
5lMWTUywGpnLcF3FKcUhLn1J8wVYeoKpb9tCb/kAevgt5I2RJuE333wDhobkvzJ/U3oPah3ioPqs
n/7uEJ11kMABTbOhonOYeCAA+0lOixe99kGUftfQTXrkfwvPAUZJ9iE0o7VqFIaqQ5YdaF6ljsxe
nkC6PJ7Lr/9cPW5d/46lSnO0ysFjdBLze6TPp4pblNA1pAszFAlOUBdhWwDV7b8dMqth7/BmyqW5
vY+029F5Q7oMYS1Dii97fI2JrQ1wR/QwykMit/3Osad+0pYbYuHzoOzWtxuisK4n+kpALDWhKNpR
R7Fk21uq1smIPt7DxmtihUzGeazH6JPZc1JMz+g2EOnVDFOzxF4pVTRt0CN1Qy/5mUhYHBkhh4Lm
3sNwOaP28a5IWPT/vN/rTSEzkyyxVDXUDJTQuiCHuLfi5M6dOEsGsG+Z9lT2D1TrdK7NyOrbdOZS
Z2dWZ4GD0RFMuS/3gk1CquTd8MlaWDxKHR/FZcLD4dSS1/5Yh7X/2D+8+80QZxr+KJ1eCEyeq7FO
DYFLJZ+RjalorhB1C8O5biw+LIMOF+bUm1WnnBAytUDL2ELDD4Tdg3vtnn+pBoa76kC4fLTfg/RB
5UAQX6OqZ9vw5sThBftcAh9+dOIrU3AEv/okIACy/FBILErtHjdqeYkfePEwYF71wMsQNa4Jd1qP
Mx/xHS6z/OWVztzoZs6ZOeflCHuEIFmF/Cn+q/uuXFtZUo6FIAq1W0+XRJDwKo0RY7KLkPGFRYqZ
vLHbaviz8HwTJijCWMl1WtTPvpzFCtMB+Xxo69g09xipfU2oroKS3XJB2QW2c3WoBl6lDPEC4mfN
pHejvmNygX0yD8bq1OkJQJvC1J00i0gEXvw0xgP8x6fyG9xnCHe40uh/Bb+aXIi6hu8557atTbnp
vJLh+sdcQElAbyleUNuO5eEMBiZ5oU7G2KHaxlwFNDz1LHGSoMGDn+d+/UKiCYZa+9+1rX/LK/WO
D6IKImswtq+Y3SH28sFpGAc6gmAJ7/u8D89712AzXQQXHn0730KQJLXfo3wl0zFYG4/edkuj6jKI
8EAdLoWd0oto3hekUIlAHV+zlyYz/dIm98PLYAcIRlnWLqAAlhhPn8aUIDMBD3klVCuN2CuOJJ5g
Fnwc1Plgs6ozbtauei/DzOs4I8biDC0bkJE/zuXLF8KFii8Td3XKyCJFshF5Zn0dfAzZoxWYTlgG
m4hpT7b49j30aXbRfp2O2C97aApEc9uPNmcAgKr5pC3jG1/WHOha2yoDzXQNMRcuuflQqtJAsiHx
ecfmKd0/rBpGv1eJv3dTcZs3J+EiqCNh93n/xHbeGMUt0wQ8Ov5cnk8rw3FZ/yXklr6naaatZ2M4
IQ42oJSkuOqL3Nv1ZXV7VoF2FFvK1Zd8j4yF2iq/1DsLdkTVQRA/HfVmAIiOdmeMqCVjVfss+BMH
iVqTrYltEfGHkdLbbtOKzlBubVmTim2KTXvURN2F4C8VXNwta4eieIoMfcKhgD3ikXKFp7n/TijD
zB3vPZVE44WW/bfnJN/QZMJx2xlnOkpPWtvNUbXXrzgKQ0WGHQHS9yAcKqMJsOEEAxezzZA7jyC2
JNTPMhO/BOrv0C47lZ0iBf1MX2U+L39xl+y9/35g0mVQz6SIdmOxmqSKRI01Pyor/5Ry9hQpyZA3
GZfQmiKQ4vixBjFo3JP4Un2EPGJSlUWe0IOiWl7Myad8SRdgXGULy6mrU+swzLXsOnYZV20pE1OI
QGYq2mhJSL70Lb6ZSEFJZwziIEPpP/mQGqwBFGQhCZsyJLLGTp0yZreSe02KIVBVBfKSPZwNjIq7
ydvZJxZgXDLC18P7FGd8iudlFHoWVTeHMJTdQXftQe0larIHrTDCFH576SGx3wJcnmjt3LRXB4rO
sNy2J3XEDcs14s3RDFaLChcnmiEtIbC314q3mKla77hBMt+BiF27KyWt2uWbzM+QW9KvxVOzY+92
yogjNWw1F0HlgnR4LDO28LLmB0Pf5W5NSjTVOKZbxxF6YNK0FQotWAhfc0Ef25DgUDO2YalnLAsG
XQwKdTDRCB46wCXVZItJ2BDe7zAeIq2Mhx9PWdjlYWeFSieZbyIXl3Mv1JtV6jA9mBWJHe9IoYuU
G4uuYgAaKtLAmm5oxWo4fa3BP9Z+wapr8auc09NRVb1/xbStY8Z24jXlVtMtceWxcn15GbvDA7bu
LZpLXgpccFuqI82JGymH/EcCIAr/IaONyutEa8YKm0I+IlRyUUaY/guZfUnD8Xfqhhn4D4REf2km
79wmMJ4heojzklPlRX844mMRuUt0qeYgRZDt19064ONKe+n6qGjwto5k/l51An5NibMKlBfXxZ14
YxI9NQP9SnHXVF6HS8Ah8FrchxTCuoBersfgJ8BWEcCupDIfgPMrt+53tWTPdggmbITZEShY9Yvm
iMDoM0a4ZmrGhl+YMWT62iz0M6XxsHP7rgjP7ikPHHNpTEQZxLdj5l42HFNTHGJuWxn4h2VwkmKs
QWFhrEs3v/h1Fl3pGzHeAlkQMK9qW8i7gimzvYIuR3JVL3coeQfPhloPYS9NbqHy2VDusW4XZAig
UQ3Lop1pP1C2He2zTxL00je2vLdaN+QrqMXjCW5WRfjTw5oBCjhjqENpX/uoxUIbBz8l8fVnhc+u
gI/1n5zNKtg/UQdEHUC1isaIkT1MGpAZMsEMwanC6Q+onXU6qbzVtqYzSEEbgGVW4IksxyDrdIA0
m718bCnqcVMQvT0+5+ewapkWJkyfR6OJCOGIaemkuFsi96aywQRSxPmcA7nyckVL3QJXkY9ea1my
pxoDYFbMbvJU/EpqDksgOPjEVdyGzTkw+cHVebce2xwD6AfbaN8ZJLJYLlmS9cUN9+6TzK5M/UtN
471VU4NPpA13LIEaMPx6l02unC/ns5eIQrZ+lFo71LzZFwcL8WgH5a0AP4iM4tMQ6JDc90nD/L5b
w1vDrYZ6EAZZa0xsN1OQtPaTSUSAX78Ejh4xguA/FXe8aU6DqcFsgGdBg21GcpWck352bW/aRxUz
QLHrWS1M2TZpuRiKhCusRNl44dYl5FzJ4IF6vI/5V6XKVvV9PPvdV16NVkDBEBgH+kITUE1OGz3n
+A0vNUuKASQPT4v82l+HmjzsEIM2uKWnHoizF22JalFZjCInk2LxSFGjqhVtJiOPxcv3mlTNDHMM
ab3p8jUvpZ+zrgGdFy90ev/m7XVbJnAgGTBPSoMSY6dEQpFvlJmqjon/50Kv36ww6I3JDKLsZpxm
pCyo6T+u/yzTM+IOw4IdddLYcbqIZjp7cOkVXaDUk3HtKr4ACe6MH+0Iw6CdKk7pR6TKBxRAKhTi
vNuIQaaRWXgBjBlyvMcOBGNf4fw34rCpM/SyjFTFzIoWk6ch4wzkM/LHE3RcpraSspoDyXthl77E
jm7OeHw8CGHVUcZYETFEOrbyxsOUXL/1tNF7to2XRaxkk1ie8Yn0nO9p/LquDvEo4Tp7+kb5XDI7
DWw8Oj02SouddGYRYtze4Y1D2pmO8OjkTTzY9c3oiQS9gs6L5XNz21nqgernRsvgs8dcC91AW4Ql
d9WQVdvmWMokRwrGqzKfKRZbcs2QaYu9DfdBwO2e4VZLkBjYvSHI5T8lMY2i+5Hy0N5O13V9pEQu
PfhP7avtzCLLPhDMBuFUergMCWrrZlUw+4UVqiJwG3bHOiYSU7yMDhxO2k+dkzJjaR2Dq/81gqXx
MTxOC1Vp/nGPDKE+hILjg40a51JFLcKz0vafzRXr5qJU9SGR9yOg63ZcX3vty4AhbidfCXAKas0M
k0DRgYIRSpCViXySbWdlk2pOlIo8/d+ZApfGqR33nbIHqicwDXRY2FpHIjd4zBZ1a0TED5gQCdnd
S9XLvcNvaYoQv3B/a/qX2nUSUXjCz2FSsX5u62erda++HuKyQjZlRKY5jeNQwRTwICEsYxGQnjcm
jhcdlFIN1u340LZqE/JLrrXlhebrAdvpNcjFtTpZ0zi6NUMSYIGiUmm115yqRUJ4tkIvv6xISLCP
iSc+wSUcQX/Uj2hmzvu5Gfx2NrgcZPa6hEaO/ivU/5peElQ532hZWPJ+aYpntkW0WCBwX5zayhYg
m2oQcg8C9VT0LQlFZTVp/5uHPlg3UeTWkTjOkoqsqvE/CDutQ6Ih804Fbc6oTFUCI7uEn6uAq7w7
rSgVDp9JyyXJxwBiV8WZAkEo+XyqzCX+to6DHMxheAiU9NJp+dQzqhP9AFXxKQ/UaOFUQ/zXheAS
z/simkVQiAY7mWyMdLdVHONJTpye7sEWQYcFG1c6sV6VjyyVsxf7ZjulSAf/uwmqko3NlwKgkAoQ
XVJ+VVOWq/iphW+85SkzlnEMEWSQvyb0ju4fccWEUo/UGd3C4BixWnQs1ewgjYJya7U18lRdOoC1
dJHv4dpEckffAik8DPa+ds2taqljfpyzxKehNjPiGevcMrEzosetIHdhUQDZ1uxHTldw/Z+Cqs0J
pbWmE9Uv+2FZWO3wOUDaX/JnrECgAyB6f/V0pvxNfBoPE/UZM3UZiM17fDgDCVcgq8YRGjwDDthp
2zLtBRrhqlsIo0Dbsg1BXO3K4QQ7G9f+BCZaOg1ZRfquCFo2rkWPLIINVS7oggkFcDH9lfWkwl9w
RPU5V7vt8qriOuGOux2tyWTB1VJgeuU3hfVxjFICcE0qkpO5unjMieaZnBhjLcnJ5mI8Majks9em
oOnNalrTwwq7y1rzoXMkBm9OI2p/Z6jXncRIky1jL6w3XQw7w10+8ZBvnKlhQ2ewDSIdIr7B4biW
Zd+gli2b0jBiTLqu5JH7iSl3N9dbqnVzQ43XxHgyqA4xBnymRSfJx+WQlp2cOuPRX9UVDuYuyDNp
Y8BtTYbqWViebsdVZ5ye6nA+gklSW8AMX2GVBCRZbayNkepBb0jcPsy1aXopYpiRJLcr5OhXxYK9
EW7sQqveNO7LBNTmn2bPWyAGrhbCZeT+h4tMA4CX97d8cJ+NAhp8nCaAN6z28JzNwgHuW9Pg/z/e
wSWcRiRmfyaDHROSA2rNkHVGMzkbz0zIlIp2G0w3IXBzYoy8ZbJWCtNokWeeEvuU0C+y/qgUu0C9
UTeVx/EwdvnwJQOBNKkmWYj3Zdb7nU4hYrppwaIh7w6LDjJ+MznSRHeMirudJ6VDWihovRBrFVzt
7TGbroEXNKR4HLEjK3y88TiftaL4bg8SzbahrDJcLitNe9cXGxGx0zMVarOKYks5dO9Q33UNQ2MK
vOv5CgpsK7Te6xwOO7d+R9WB2RBQckdr4sQTnwlwha7tA9F4R7+lfwCsw6os9iQJkneOBQPtBeeD
Wv2IuKgdkcQ1SvTmusD6VerY2dexYBGVeFM6t315XkUfnrNuoF4SJvLVGmC2qw0SJUyRexVlgNsJ
ETCnxFO188ZGtOyIWnbcknGmEDOv1CK+53q6lt5h10APcAY9ZiWHLxJ6na05J/Svd5r51B+4/6BC
fbGHi6zfNVDAnaeT8T+JsKww2fKRJaMxXLPHGGbORU14RkjonmEPWQ1hl5zf2z5daj8ZBdW0tvMh
fzOKVVtRK+gbufMQy5dP0PJZJDGtGPkn3cVptatnvGOB9158RmeGaYDlF9YU+WV7jWzs2cYp4vnQ
myzRXok81ss5YpdAgG9+u6c5QOsZ9A4UlsX+kAaSvxDgV1TcHnhdVWe0aNB82NwPdnSf/ZfQ/GtZ
iEMrNVoBj0r6t/zW0EL8/NzUNl/rbYx84FxoruZOephiHW9a/7NBlv2G5msSfm995/zNUwG5FMAP
Oxn67jx0tSd7aQX87wDuL84t0038inlRIP0EZokZHFRRNZHbX9dLx2IfAIgSToV+8DOAGasExlwh
KB8dwb560aJQdZGDyQ1cX6LGr4RitFfEAMBnek/25OJ7nzE0JboaTY00lNEhq8kvL1UYu0Woa239
vKA7bUZwgHPrEjMySooVst+5Xu2/Y19uWT4Jh4pHNQ7dl27ApeJpEK5nPyT3/Yp5kpc3VNE4JKzP
tnsGO4GOWoguzVE96JxAJ+F1aHlNMEWaS/22CvxBObmHa62PSCllYe6aveHfKMTtoE1HeTlvuRxe
nxT5XuCbcvMg62q9oN5h/T0PzW/0gGE/XngGkkGYqNTC8zrqq4naRJCG7tibrlEjIcQY5o+uGAIX
fcDfe2XJx02JJh4+x8xtVBCCL/H+2oBFzO0BXG+cIbm/0S4yednVsFzyY6ic7lMuL2z+LYS0NqeZ
QvT6jdIXMj//3mE0viUgRLVx1PIQ2bf/v/XqsgeUAl8lP/fWdpmqicgQQVM1AvB9DQsRKt5Jf1DJ
xeN+lc/Ay0z0006YC4rw0wjs7336gCDSlPU7Cx7ngXLylbOJ0P0+CDBQSUOk/Agc7NGGNK3k1GHc
ETMf0w8lUEUPbaFPe6vlxV8hY/1UsRr/EBO3uX7Ph5m5TsUZwnaqVxFvMeKgmnQPuQUws7WVcViB
d6P4NlclW9MAjsKHVlou+SmHB6PDtRbg/23SO2LAC4OksLleEPfupBhnY4K71EPBEo3bpa32NMMY
IEHmfEmKcucn9VxsPTqTQuvX2/DYTHpDOrvDdrl1O3dge2svos03HB9uETHeYC1aKOqPlnOBApx6
EzJpBKfq6z7cmmBjaj40/t8do+ix+y9KIQsGNt2Vx7svKXN8LFcUPcOcjGzAfb98pPdi2BVhdx2C
m/TGeAodZCCiNLdCckz/HpsuP3fOMt/ViFoA16Kc2fA18vZ+yU4tSR/pO3cWWdIRQEJQf2eyanH7
5XRjf3/qcQRj34V1ciQGrHL79eylC+i9hN5KqtjSLpiNaf8+NYk1XypunbzKHVP4xqdVYK+5ErGS
+3fQKk7Fp6CPP5TGiPzBW3e5fS8x/ZDAArnxynJuEgBM7qFQcjMt5cZwo2dVCnIsLom4KRoRnf63
y9GNHOG2JMzORO67k0YHdk1qJqE5+OxGubiOiB0LLQAgDG5k/EczN2/YOEWFn4ldSlxU/5QzMiHC
JayPE2+F82Lu4oUqnlQLaGhuZ5HqvpaQJrHHpc9LhXeIRLbUDWTLKVAMOCGEO1rNKKW3BpNfzyM1
aK5gtN7sRGr5PhmwbRmkGzvu9hlO+coUCRA/Naqp8iA9Y34ecckOdL+qS6+u4tlSnkHah66cj+8S
AJd+/MljO5QiJBh+Ap7we3T4kwbBoohmbboGIuah/qJBzIYintl49qQSeT/2XRqKs1ldNn/FnQ+W
E006MYLsvZspa9DrR9A6kHMQSSZ/WipMUrx6rMzAHvJjqkzISutuTFScWhZhOACkU4rurx7IBuI0
kqE0WhdUmBdSOWQt9kFtvXlMzBlwpA/6w9kdEN6WZzmoBwxF2Ce15cZA+VQF5FibK7JDSTc0kCFx
cs77XQm1M0DJmqPpYcPUPwhk2ougCOo8INtomHHvYeRLFvSU4VjJlf8wWP/tDVCfwLSaYP/Wo7O4
ea9zzhyA0EBvtc2cNQdQLNHep55KwWpfKQewX/EXkdi7tnbwq6KlQ9DcSEUsuHYdccoQs8aM6rd9
+h5/16sA0rSFA+LTcqOfO2fbkZuyaA03HZJEH0lKhn7pTRhFonqcCNCrjPjdWuCaHcPHLN4DBXgz
3tn8spdi6mEYibILkIiStAPPveYWUCllL4O0rULqFUpRykKn8hJ4vnEd0WzlUBKBjSLevBnNKrpx
TfCzyVR+JI/nVyP/I642isUAACClEb5z/4sBkVm7Y/P9+Q6mSYLv0XoHht1U8Y/XIF7KNN8SNr+K
/18OdRzkug0fmJnVfkcfQiu7Xsb9xjlHreNDrTY6N7WY62dcgScRYnKfzLrRDobwPokYpV8mnsgc
DtGsx+TlJHRbG5zVKBmBy+rQntsuEXvuGzlpEQ+ztIayzGEWAfnocBaPruUo9S8MBURyJKq8Je1T
2DRcxgaP4EmS7w+0e9XN2ER9gYLZ0V8ujx0DXDIA5Nr6PmqhP7/kh1OaWPac00hXFMHxRwkRDe+1
2vtbBMJUik1XCh7FI5D+Q8hVRQk8pXjbNSp1qmO9bi15AnPrmBQRlfBB24dpHk3WwEQdkQTI/ioz
qXizxAr/5au3mbGlPxFHDxZM/wnQuaZbNl7YW+inZ7esdZP5Cuy3V+YH3yXqWyM0+Cme1KtKD3LQ
UlmGiz6+omh+Q53+zcG1y1aDyMq19wYrOX+jvF3/QWbwP7p89eIndVEu/PYkVRqLxzT/KiHQmVyo
sy49fzp2rQ9NnQti+bqJ8DgWkexkS1XYL2hP3fMCwv6smK3xHQApLLuYSgafsxwteFxQJ7aBuBwV
1jOT3XrhRhZBGQSGj2plTklKPbTM4ByOKYFZfLTlIF6vIYca9QdmUHC1Ou/4qG0fg2ByOH0XRAlh
uQrYHzxd8eQHJT346yazosY9SPbqBJkts61rG2qsVdItf2CuQPoB/v1CgF+r3/UNg62CJvkia1Ay
0EtGTU2GeyCyp1yWJFFXMNiqtPK60VqkFRZ1nTk8R8IIdGKTFqFh2DxWLHdjFSbLo5SxsPEGVuy6
cDlb5JdOLGu2Ab608dy3w1IzQ0hA/bGxA+yvXkYX8Z6JuIKYQvK8a8qomCX0OUsnPMB29z5rC3Bk
Eybjn8bm2XYpEMthEpUvEmYmhsm5sTSGgnidZBWZ8xbLZNVPhKX2vkVWulPY8X37kA1bbKBLlG61
P3Zy1FO445oX87QrRskHyKEuNnWjtHv5HB1K2MDCP44KHRXXLwlss2EbBRr4ygJylJKfbmx2p8gN
mk/K5Br8vooVLyGiqt77Ha164QwZhffA6Rv7Xq31R3uOQ7wbS3wiX8TY4Wy69GggnKhPXKqIJ1Xv
SDJWB7YxG8UIFXJ3c5w6S1D/v026pJYza9gxw/5hqrU0jC9zspm0vLxD9zZdT7hGVhmcf1UUCEOr
i8UWrMPQhREXvIX1nDeWbX15zopxeF41t+p5dVChxy9WO03MS70U77Rl/MJNmARY87nyp8HLiYP3
96qb1lPEttRbGn3UPbQfQgD6x1jvS04ZapDhgPn6Nhd2sCdGqTWOhA0PU/ObFV+g4i9wFNFhRM73
ds2+BM+9t6Hgf1F6zmBgmw2z9U4sD6QaRwhzjuucvHnKTQ1uxeaZxyLiRVYanZsTBhZ4igljFN9o
E7by43nf6AsotwlZTMGhxjuSRchU9zm+Zp1YP7WfPWWC34bLi2y3ZZ6iGeSge0BvYHrTBJhh70uE
XYkHayG8+KTHsirfn6+VSnSEFsNhzDeXlGWL2nMAazpa37QOZgfWRtqKICm0s14stlZy8lr4aeZ1
+dvkiXzhCcwhkGECfnr1fnOHt+xUGhdVxAC0+uBNKHDMGKbCZQaSqESTDZkorYEaFXIQVxTU420E
IGLJLvMghGibTi1+oITN36/y5pJNUXVGOw0Q70+f6qUJUNiLJjQ3iuSXxfkcZoofjxJDcali+8yy
UhvmB/nKVsMdgEMWBWGUG/fkZwvkKVPXSRQwx6uj9MjXZYQxpMVMydiP12ZO95d6xLwCkWLa2pb+
C4RY8+G40wvLpp87ecGmt/l/FDGKaLw6g9mAcqFnPooIbSZi2M75Qpy2hp92Ptfe1pOvVRokWgRr
7LFN4kfPA131tsanE9F9LAFlTw16slJoQjdpWA7eSd02BaxQDMqA4b92KsFmERJ0+AtY71lH6S8H
qKCa17lkGBa2wTciP1+6uubRtDRfaZG76357C8khyR9Ang1sgueN5vCseEfxcy5PsviTgfROVOZt
q0b0vat4x9eHhlYziSrqFC4QbuFOvc5Ic+RvreBbxbZMFr7qO2kiFMZ+LcTprQldUAFFrFmmnB7Z
0EpacUUy99TYEB+xPh9v2WeVnk9fw39kfvW2Cy3Of9YJ0Z0Wl7oxWUzBZbf5973CmqS82cyZCaoH
/9k/y9KiE34zvV58gB/Cu7mxImgflWXdyKWyZ7CHh65AGydxXQ1GMwP5en1JwCzFVlAuyN5qlUiB
swHdyIuJmXMEioDwXh7EVyEwczJMQF+8zFzmOBv8+KqW8oryBPlka7pnLQ3RElOpVcIsnqQ2mA9Q
kdK8P8aiPW/Rpp59So4eB+2P2GHCIf1w2VFybcpLWq6cAJPX1kb9NiaLOtecSDI4U4pPAzKXOPrp
75Ni6vKybrhIoKTL8hKiJnIgZ3QNnajGJ4TM8MRfPKiP59Rt99kKv4cezlYu79JuGkyKLWTlZawI
hjmQ2UceJKiVBLY4z06Oo3ACBpbY4RDrTk961eOTVQOvcrUej2QBlpUMdeV8qs16VGlNtzEBAkZa
sAPm5A5av6uiYCxxEgGAU1LQk+C9Eg7x7f/FzgczbZDXirG+KcUlJLhNHdM6A6wcVxUvn5t+yoqO
D+oSfe7Lzfumo4nB1A3uHedpKjTS7cParbDXBwP9XJbmMFkit61owCKv9Z0raJEnNHmykEwFGkB4
+GnqB1madDh/2NMbG/vP/zVATdSX+JTCK9cTavRdFWF48Lyr2ueuCBwiBD2+4nnttShLdj+1Rwzh
A5H/wboZpd4ByMUpJFdkfcS/lsIO2W/gthLYmo7S4JER4/J5WECP8NoYnfqgm5bhnc1A4OcEWmxn
F2CiHHNi1bGIYdz5q3SqM+HkC6erfzigmDNfq5M+BhIkmz/xe8q11MoIqe/Frl9RpBagyL9MfRN+
lBl/OSCU59L3IOWFl5Fi1f71QvdzL3TyNqJaLpxcyqHW5EeCG8p9hgzMau3YlfYFspYtrmsIP0w9
35XpEyVPpeNtpM23MM11qF38qA1nJKoPZhoSQdPZSOnk0+YhS5bAWvYgY6T8TNkjrD1V5xWmse36
Z9Ah7H11CNyzvUxbt2VftMuGISznRqHYzNquhbgr/t8VvKdPNhEqvz6eJv/CWRjiI5yHPAhW4ctH
i1GL41IDKsdkCEBaqJyKVl+B3WqByHRau48HRaUXY6Pvr+9+v1Fb+P/GH+el2De5mz02zk3hJ7hj
QbMyOZz7RgTpQ2lkifC6Ijkns2R8uCG0tFWhVMbS2UZp3ALp2SkqIwNz533pesQHHu99OkUmcsO4
4a3MjsjVmFvT0W/IgRE/v7xI0ua3tvA1+dM660tByRUPTH83cD5zWnlEWplDvaSKxvKBjyWRXjFI
IZJsEqB6yF2sLUwQLpXLYkW9e7SiSeYsEA2fKZildhWskqJ13pU1g1ubO7tGH3V20y2lisPjHsRG
yJko1CgY4Fk2BzmJr7bs6OfhBMw2QnIA0RNRtsmrIvA2HE7nVf5bNQNBdJ8auQ2nIpUJPSCIvxdp
GtqS9hitAljt4oh2hdnByEga6FVDs8HOupEKGSd9Oi95TfO2W3jEJWVvO76BeIXQpsFnBH1Xg/G6
icbBRHxeilu6XUCWz9llRpN+58dtmWhD0nKrX65qMWzAo57Uu9S+O8ohsCF/zMHWNu/Y9JuMbq0f
LEaD0ZdzUvG8QzN7rzTUbVWd32qeq7y277sBZozxuF1YRnzmLgp1DiJA1e5hLNS3x2z34FIsYGhC
qEDSTaKDBT/8ykBcufKg8flP9aK/KP3MxScTOo7P9ksnt3O3SqBAqxP3/eEYK4+yVPJk424eJTBH
yU+5k7hEPJWSupQp4b9GGWOOiLCaED2xc0o2sn9xlEbRxd7Enlb5uk63N4/KOP+/Gy3+1iwthDuZ
iIUsdkVEZEnPmtEN5tkHDIhF3Vkf5MlZnblx+G+TzyQimVjLMAWYlesgW6f1D38wU8REX+21G1ju
T4O4t+IQDK4Po44N6DWrYs0uxgsf6t8TYRoRmQGrEg3iHp/SheebNwKx5jyRwEbEHhSrr0Eqp9Ni
7kNyFmtVMgR+rHeD1l3c1cC77D2wZrdWEngSBd8amFEDzo8Wh6F2RnivakwlTp9bBtLmRm6+WHEv
r46hBdq86E1jMiLRWJBW5kb+iVWkVG2nvPKxFBr5T3ZyVF2tuD0CooD5cKFE1yxcAvdjOzWyEBVk
EAQIQ2eF3eVvCojtxgW44JfrEKo/+ak0wfFp4at4M8TBe5T1Eoi8OSH40kcrQTwX4oJMXMwfJ02R
+iaC68j4J/Vjd1wmeeiionIrMnVP7Q2OvqhLQlm079Cmm0dnN/iAcWTelFnjRm0SnDvuDuJrkP8+
9BDetE1nQtsZWBmdwY2AWVfWTIVRAa0GkIRBFEIVTISXbnqW4Yg8OFC4e/qP9/w6FD+a2rptUpWb
bOAEHJvZIPywPmx9P7nNDBrdIzIzUqCAc1Xl/SASlHoXhjgxl2kLYUAFsys6W9sNyMErDdwQbDrc
oXAL38h8TGP6hmP8ufSOhqzUm+KCD6i2qiXXkne94W0pJsJQ+ZLu8kuJOqs4l8Uj5BRiWUTXqYUp
ueAIEh6jIawIh/7+NxMoIZveNkoTa2b3LW45fx5hA1omJcDub/WwWdsP8mIU8GX8JpLV0kALzn1S
OeW8X40NaH5rPOSUf+6nsdTdqhKbIMzKgqGEZA4Tay0Gs4VgYP+UW38VR0dBxFiOnNixCD2gOFBO
F9SeITAK4Nxq5ayegGAQ/YPNzXjznBEjmncNbC85w1uur8Ds2yVKrokKJbmbEzpQc5h8X72ldqBL
SX1OhhtyVVUznCGoxQr2BeTN0aOJOpZ5oTQMwYmV8zx6y1dFs1uNtst1oLmrTlJo6yqk6CB9SNWQ
4VFAY8Ga+BVkrSnIUv/7tOejg/mMcxLN7uWerNWu7VCiO5zkoWbalJAM3ypX/lWvdacbOGuJ2HoM
vPXL/e6Qao/GztdrQexKEQ/pPJ4BB4yLhp+INsx97pEUrCrOduXGSePCwOb771FE/R2a3ZxMDj5h
z7MqQOsLCq6BXvDcI9e713e9cyP+GO/8B3j+Wf1H40E4CpvjHnTIu0/zssfdJR2TT4AnBBOaKmnW
x04X8FB+Ofz1mEuuljvmNjbczNweZNbAWyrXcdt21AFAC2cOrRIRg/WmL/PkNXTFx83OgzhEi8TO
t0HV2RjlQeG8lPlgKUuidDdvpE3hjHVdPo0ebdFHwfHcCSye7PL1WnOGKl32Itcqj2uCcOc/pr1U
aTB7zao8955hpUEFtjHPQyJksnOEBpb8tQdiuzb3uvpAN7BzAnovrkhUFnR7dnEXrtKHeypFm/8N
7MXJU6tOx0LV951WocK4swb1kg+9MlKVeBlPQ1iC+yV6ix+TaGy7eSR8Km3mK3BcpiRjbbx+I2cS
InogU1kDLFC40PoK0LRLbqXSn27h0AMD/Xu5ENMYfGAdVZ0KLmTtCXjE1VN/zm39x1qphRPHF+sn
6JsdVHVps3FWa6AECr20kkf1eHvYuybSz1HSvtnAZpun0TroTfBMXk9CZSmBEW4qKgmmYnmORUrM
Hty7yL8QoXN/QjCU4uaJR3jR9qbXaTXOP0T8FoPtYsq5WbSxEcRJ/wg5syEV5p8aq/v79zXa56ka
950ws00XWZOP4ey6z215Wj/Ht0Gl8SrYOws0UDR0SLJZwi6q1ngUGPfoMWyXOBW3qyFC15BgnT2p
+hlbKa9a1OLzfx1JG5BhB1YNkbYV5rWZgo7Wh0VqU6to6UNCM+lXc1XweBfqGRq+0vtKpSnW2egz
Ahdq1fOf1X+U5Czm/4Yriep8s25NXJuDFkZegyOC2RR/qu9Kdt4XufyIlmb/nBVHaqkfL0heYWqu
EyIk3oKV1IrcqbnC+AcYl91ZU/klcnDh/4vBBufO8SDW08NebaDI+P+xr5gBD16a922mI8Z735o2
caxm0a5U24hExGd5Qi2CcHK+OWa1n5TgzcEitnZSFXg38Uuun55IxxoB2Bt7VUCNaW/XIuZO7SJk
cnt4cN3M2FI8ks6rVEJo6u8NMalxzzkLG4js7dNEEEmZ8B6W8qTAQiMqVrvSPSM1YvaNQ9cx2D3C
sok2kfH8qB7HY5GMw0RaqMv3J0MiPrO73x5+KS/bEDMShIZ7jdSJ6XAttYL5vCwl2ya4w1RWKwa9
BQA0HXdNUMOzF3Lxd9YlKS7F3HP5xzjINDAfp3T4CzCRNlkoQn5IRCQ6vWXE8Mife6ti846cywKZ
W6ZWBOUMyLboeiLN5FwR9I7DJQgafiwkXa/655l1VFbT9F8LKiQPRp2F9MWhRuewPsIx+f20VlGE
FFAsVvyjYkCr+u4JtBnc6tx+VF0GBW1VjmbY6eZ6X4hjXNEgUi4EKKnXQ/ZuVDfYtnaZH3ksxC6l
8/kzjlKw5sf5I7zjP9svXFPVxptKZQLRstUl5j5Ty9DeLTxzySOS2e1ALrD3xyOuH7SfjlzkzkA/
3WQlIxNPs574PrsgJuvzIZyRHVQtdqMVCjjhhHe+B5U4QCjucr54pmwhYKvreB/T8nRl/Y29K/rq
+t3Wo8j8CGLN4pt+/5r1bOayxdlnvt2xZ/39ZM/OiO8uiateqiDLHo+BoHDviYCqg3TehGYbDt8H
9gnyF92Fqy79Y6fq/vV/cFV6EYghtmNylVT2Ixbmd2V7qExB8GkrmYiHmo3XtQTmWxbsgymSGLxz
qXsJ3i5QYULCj5rQKsNv3H/RBAM22CD+bQ7qK4Oe2lfayl9H2g6/52OUUjErheIxIdL05v3qf1fl
QNQpiNtjaUnnYQBm1h0NbkpbRbX1MscW9FepO2GtIVxUdY6HM3lUQ0G/QOlnGPhrf7C357eHG6ZQ
/sL2KPYw45GqXZXNtOi2+WxhPS2l054uc5QHljgJnP8KaEvShEYOBIsWpmZavI0nBStp0MENfAkx
xl0PWiEXnLb9UHb4IteOTeyS+HvSIkUrLdpXLnUGM4R8elekZjbiQ8ns5HEv3zG10ttf8+hIC8pY
XDEEfJHW+WbTt8n0xKOg4VDvgv0eNfJdTJ9Kw7DlA0kodkZyfZEfWlE3y0YW+Bdq7XWOAPO2afuk
dfy6z2XcVWzLh6LObkNf0Yt0IuvifsfPqYjdoUPeAobWJWMwVeDtIu+08Xhwv8dssMv/+oTiPEZc
TL+UTEWHG86pa4Ps1FIUkxFaUzr0f4388Hn0/y3dgo0iMAlJv1e8Nr2CvxtbgbJ6rsr+0Ofn6O0h
MEJzOZdcFR/5G71xeaXVWcqmRpPQ0af98SnW2mSGBU/Pz2eSEbwIJ0clqYNVoH4XcDI8ENHb+l4f
uB9ANGMXFCPsGLxHjfMmhek0dagyZ+F/7cfkeaRdr8+sXziU4F/+1Sp3VMcMzDPAgPjGTc6DA7+C
xkm3qx283uy/S//qe8LVw/ov9/RGtoHl+G3XrjMqs9sHQ17D29kdlx2xFfuPvF6yZmTQMFlz3MWH
3WHtm14nlioX8XWpddb+7LM6wxLaq/zJ8fcqFhZfa+I9/yKKbFZMPLWlnZnFbFK2YTnZDlfr7mT1
/HPFKZA30ImC+6O48I2RatITjn7Ho0K8OaMm6eF6xRs5iAroCZSpyt27n2TKOLH4ziZAe+ugH4ef
4jNwEHIbs4wd3DIsvQoZM3a7/QBB8uWFJ0I/lbxz7yPmAcmUwk1wPJ2KMUyjD97NR4DxjnVK7fnp
K3clQ81C+TrlE7Co1+mHFlu2ScyDD1aIrb+KS9K+117IzEf91LO018gPJO5umCy+Zjy8QVRomCNw
6rbs02nY2FBhUndT4dFMHRHnNEHIdwJfrzhFLkiXOsGavN4jV6fffe8cTYRRl06V1H6IgnC/kq/v
fgRpfyg/P3WrjMO0fWxaBSWvsTnx+ssvPLsGSnT5WMPwFiID3P5mtCr0bhQaMN8wWUqfZeeChUma
bHbQgUtUiE2Mkrk3fjGPgC8jvR/sMVzhFnDFX9vHO+uo7PjPDU2Wcefor/3re7g7EQs5O+ApbKrQ
q+EpDZyvxOTdQJv2tM36zVKAql6WQBInS3kiZc73Tckm0V/4P5IoiEqppIWd0kKhaxhrJUhxvzQA
X+aoxDDaxoEH5jL0/vuOC5fDkUdOCkfLWPDt+vnDGDLJ2wNr4t+5b66JjUO6Fz1Hy7Jpmaos4hKP
/iIHFPJrGYFYNrhMJPJL4BhxFnYTBVf+CtFzFcutLRfIZe1HhPBS7/z5nP7L+ujMxmsCQEJCw5ai
SXyUNbdG6pWWKJSp7OLruUwFJgV5fSxkMREtewyPo5+eOs9Tldd+yCAawophT1EK/Ah9/kjFRnPY
cp36ImeXX2sYlCPhL40yipioJ+8pmsVH50sxQRz5+X8/t6L6aZkwjQDuW0QvZd1VYyB0bZdRJ0th
Jvk0uZ9KAhjU5fD7GyOAgmZAEa1e8zG7Q7OyxooTDi7F4bVEGYi1SkC3MlmYVR4KDpUS0P06YG8j
Ogr2662XduUnot+qosc1eB/SzAzpu3vu9IbB4yFSnQUFa77a47sCdsKiGma30+gahC23aWpIYND4
dJhH3ZpGOo9fw+Jo4XmisyuvYLgvrYVXMzMuFRaleynmyTmFn+l/8Cnlu178k2IoFgUKSfgZp/Ng
r3UGPCIr/OnCMdxbehTOYvivxlrp2n8eHk4pIgQYXPDudqSa6Zin8fRtK210cjVSthVRvCDY9QXw
ec5XwWzHX1+Z3EGIAQt/lGAurhSFUlf0O+E+JrinlVHELgMZLmb/jXiMZiFGGQ3NZh9b6o88R2JX
dNWhBcBmDdr7QgIcN5BpKtT3WyyFfkB9FG+l1RmvY0Gep7ctb7CsF/T1ZUfUMtRjZMQpmP1ffCJX
uBZGX/igPXYXv+Xl32Yw9WQQ3Gx8S+0ebL642RG+dqw3kYWjiJHT/fpVBhYe6gSKulvpMceYTAVe
I5zo++ISimh4/rjJVUS/IX1jo2E2MdIJ2hAUMPvMsUBMw5Ht5bnx2KuZEn5wWOLBqifhHbujMnOo
trejBooxCQ2xLBCikiMJQwwi98VdCnGjSuIFHEuV3dIwCa7W5FIiLdG0bQz/l43tETtPsH/5tF4s
rqTOX4ZZxP4fqPiSl8vLFvLo6OKlVPbBUgGCtIdz9ZpGNYnc/gqDfk7y9XEeGFSSXoo+omFS9aUF
j4QPLwtfN2F4hR0upjo87l7HO5jyNzp3QAmx9gKthKGK7Hv9iwSYiE1CE1WzLb2Igej3RDMrgiHl
j2hirrT3MpQ/MQ/7RAf+0t2Ip5qjwUoQ5UdZv+rm5S+u04Ozhphdgt+tGX4V8gsMpegmj+ou4SNu
1KrIS8rMGBthr71bWbKtv86Io5G2Y4ws3jR17Y0AGvD6D0FsQC0BYkoEyXo/nwXtp9iyzyDANWYq
cuUpnS+0wlVEZ/oB0weorbuJ6zrGoMa4GZ0ZU8N4N/puRRXHdtQ8ZuBGos/K4CRS0X5fdhauiJ1a
i5ln7Ec/3kWN2IXYdZ/QirbDfWsDMlDLOr3INgFBk/OXf+7Ha4x0XItizc3YLeI1IMtkT+j28L3Z
dKr5nV7Lw8g8R+5/C/sVbQWF1mu/v3BjIUK9SRm3yB4sh9yryfOquoC9nK3p+rFP5mjyv8+iLHli
tdoIkAIbm7uqrtJzwr8+zdO9C64AJavZ3977DW0fg8YaNqZ0hx4m0JikCyw8432BwGUNy4NrcXKu
Nac7VPLR0cYD9v708rZR5rCAXA7pXsvjx4wpADHWHJnBOZFIb1KlIWDKGUeAOoRcYflWmVUjwFiG
qQDUBhZgRx8ImBmiixGSWdxexZbOVP9z1q9A/PCw1Q488tpSvGyT3Wq+4iqQnW8EGGCcfYUzPXcQ
ci7YbnukZ5nbMaU55bo+DsoOhhuiwE1MG4YO7sXExHQMcpuNPKk2XBC/muXj3iAsjbSgT4jJBQqh
PJuIToh+VBOZ2GJbOPjY04om+zbbPCLmn7SbVjv3D5Rlv4g8IFyIxHoH4BlbJrrElRphtDpaywH5
v+18P16BSyjls0zRMhcXcuhsSXY1JItpWr26yXLziyJ0W0w5SEb6d1+HMWcKstI0xvItr2D/MhRJ
O8avVdRm1mLU0NXh5tPh+7694OqsFr1iq5Iw3TOv1orcJ3/9OYVk+A+7PqJY4cCZUMvQlE5F382R
3oQjZDmfAsovrmAmsVSFFQxUG9b+l2yB9IfjF8IKs5dV/rc6hQuTQpZCg7UC9x1y+wqXMEPCcWRk
phcqtZn6GJtHC1RFVwfVr5hV02J+4OX/ezaTkY0ktydrBgByuB9mcZcjyrLXik254ZvOVIsG35Wp
Oz3hI6DYdy6quEbbu8cjM+a4gTl0dBwadumaS/s/ebrFcoIxpxA8nYcMiuvq6EbFRzhbNhyv25G1
ZwZ4mQho2ZcVnBx03IhdPzrsiHtGkWXPmRDR/yhvKerGkLkzXdWsIXRahgFwaOE8Hm1zpvubLjDQ
/8TIR0H7ROAaUeNNZTU3EGOXr3jnL379e3XkLAif+o6c0x0eE3FZhLTFnIxez7kKVrS0xCg0t4xL
N7yXN20RvsUjwTqKt8SEuBcfaCaLj8btjcEwYgBFWJn4MgyjSuqnrD25KwfHhyzhUIclhUKWtO+u
kft37DQPlBRHqVNffpS0KGZ8O6PT2rdWdWeuVBBBzNEWz5aJlH+F20sCmlw3N6NJSvqYeD8GF1ye
RdfB/QwrDpdtXvKD73PN7FrXiCq9KXEcV/9CC3mjsCR6VW0D4fGSAdvBIhIhpUMdY8oFN5btQ+xs
8qgpGbCbnVKMF1dzpsTAa1oPrYAMqhQz5n7by0oXPAd17eOG69fRM39FuUehez+0RE4+Es9iJMU9
aNcnN50B7kHhrtieurLVbBzZugOjTgKr2iwF00P0qXVHJxVxCfhaPrEbFo99Wt5pFwvQ39Brg/ua
GmxxvFpArYxJ2nd0okBCn6m64LbtM+p0OufCp9y4C2q17WxzyuNeuOOlxZWojq+8nTJSHUvERrYz
rDR0ZfE6tlbzffy7cghu1ZmGcW2QL7AVb/nKw2lzpZxbTCj0QHhiq8h9e+0/2GU1r23AEG61e9W+
ECLco2cQgdeQ3X8BAULFma76CA725iLclzswdCvO0IKZt+1KdmgHWU1mn3CRqa7V0sgGx+nrlQjl
/GZZrT0g5lCXLe+2dBB9lBQwo/BRptupZuKpzJQxUWhDMx0OFDEqWPLg5qMUNvVqqHrJaWW1Kjd8
tEiOXFf2JMWNnIi9OgrHSaB84A35CvZUWgv5143Wm1dBD5NJC+wiKnvmUxHpiGoLGWot9jF+Wko9
hg1o7liEF3V5viFac0geimZPFR6Wtq7Obd/TLCmgM+CExtcjoLmwq3BGNocbtYZ5D8Sv1nSb+HZy
nKanswg/0M6HSCxKAEY4d9EnEw/niZc829TrZ+XnDTZFWuL9AWzksd+DYHBfT+6Xyu/mKLAyvEz7
nebT8T3i6m4CtyNZJik2QzIFKYnUUlwemQCdycolEg7Q19MsTvnDmW4LOwS0qXF8kf9X5QfrkRQ+
M02VzqxWjwvI3OVaeMJFq9y9d5R0A8cv6CBJvav6ICSaR2PbFMtpZWHHM05QgvsxfqHrAYadYOp/
q/q+2MdoQcIss0mwg9aTJA4XF02f6fYcvFpfNrxjZ1VryuasldQhdD3LgfRCb+0gA4vS78Hxz+O2
tLoobEn5eR2XqQcDk8U6P2NvdMWxBNNnZ8b162JB/ehYf6FsLOZQuwtVqGmGf7UXIDQk+TnWsjmw
jbj9ymqxPEQGO2DxzEFAAqCLcmh13CWMaq2I6YzS/V+5xUD+K96gmM02He1S9AWj0FO6NstdXknP
Rh9fhulTS7rp5jgVh2WNN99iV/LX+QZRpQyEP83zlpaMCT8ap4emwsuMzMFPECH4rDnp/hDcNvhW
+gwyw81j9LX9q4Iv9Av+tZVt5DlAzCtfzBcOb1nFqX4DRBFxDtcB2C05F5WRJmZOz2iW8LunKg6K
LptF4WRiJimtxO5V5mUdhNZKUnF5WlUWj2NwJ01Oasr+YKFn3079BX07tKTv2qg8KfQRGQbFDMy6
mfD41ZjCXS5LyDO/KWPnSQRNkWW+gLNWx7NtkRJ+MlFZJj2GJirP+0iEjobPYjVBQ5fRq0/s25GM
Ua8KZmRm7gtlmtyTez2F2Ou80Z2u0GsU8p38RF9X1cNmxQVfiztydfHRTgPCRl/zPXTyyobnHcgY
g6ioPI5cVJJjOJsCVLWyLATZZh3KWaaRN3cwd/QYAB+XB6ISrxo0/MsWXJvJmBLa4sZ0osKQDVIN
jfheV5Rhn/0Vfl/EIhcJxHuF4v/dQ6zO3mmCBwX8nUKT0tG1A5uCO+3Bvjy5qzdKEqOOvBt3lRMc
t8huHfVUJ9I8rvalG/cN2cNS7g2cmJbmiQy1I9dDuqo7wVMbv11MZtlF1fUPNIBWQHmkYur45hoj
aZRNwI5uB9Ol+v7ntQhPRp5rqAyd95NfuqaYss0RHeHlb3Jy7GivRJtGQorkX2PJk5EYa5Rbx/j0
6DjxBR7kmVqbSUxeg5mhqe6doQIV91EduzfUAX9UiAHKeLXyaeWgJJ8HII5szsHaPbUuPoDdzxzC
Xz+U3dpYY3l1cuQc1F0VZZZeQVkTPYTn3Vzf+tUDI0U7NtAmiBIdWsq1jtdqISnj8quUQjnzHI84
mk3CLQFzeitFAJgITl966V0+PbB0xpJb4nm5TWbnBSQCLQ9Oa+pyKTD6voAPSUspEJxHr7Vi02uD
LD550DUuSPR8z9lJFFp/9VwR1V6rZPo1N6i5CGtKvFVeET8Rn/TyOa8R9Q4bXLdl2/WvZujqkz9p
42btOz/fHaWa3Jae6kRql1PmgXxWEcOZC365ZeOYcEtFF2BbnRNZwQI77g8AvQ19hqIRMAU5znYA
yCar93XstKU5WPkEIQ6Y2N5szn0VqZbKN8rkWaqadWE0V0VeBcD+D35cvAbWRAU+i0/vem7q29/G
dFc+VRAkVerFo7xsdfhYigui7IkK4HbA9GPQMtVC7G4XomO3mcNMa6sLheu2tgIwYARS438PHsy+
GuS9psGq+lAGl8oze09nd0c4Ts5mp8dLoDSmdyTTqhhNuWDihwn/reilRCMwaDSt25oTOLwf89oE
VnZimuCO/q9+1HLaKRYeYCrdZe1gdM32MjbVQSP+JS1P0aku+CiSFfGf5SNkm497Q17adxn9VZny
zRiSUD8wDXe82MpK3b+7WJ7fYJGWReh7WYPfWMKAzH0nWgx+36kyvebMryImOuU1GKzeuEPaElrn
gt5zjdlaYl5QO+V6absMgEPrOR1P/6adGgzjmanVFTKpUQEFu1RY0iddAHWqQ+5oOnXR7nSBkNAV
cwLuk8TucIrp7dPZs4e2NR4gOTvoeYEZ60x/l4JzTmUT2YgCfSE0joLhfTZ+B4FJ4RZPNzBg9b/t
ZFEJYivK14Y25WfB5Y95qRviITsY4qkQ0z2YqeeMF97uHtFDAUT+rpb/b7idyEGJK435+G9v4DHW
ebrGi9x9Juu1lnHpGOhhsAVkMVNihNljNQw0SMEe435ug1OjUPfgo3OZxFoi+gvBy4EaejBWttUl
uofzd2neDfeNJmkx5jP0NfQEZkHRlP6HpVVi6+5d6cCAVXRkG7zPg3a66jsCs+cRjspsNldkA0yr
B6CpBNDsoR6biNQF+6s4/ekG9c8R/zDX8F4oS6gQkjWrsxxSsSEI/JcqF7XC4U4jHgzGjf9EpF8t
xHX9lDrOUHCHa2aSuAuYMeExXxfRHQQXSOewagP6L3wxcp+lIJxFanw31MduLbyYXNzYdUSk39Es
b0NPRo4IBY4i/P5Y4CMItueI5gjlsw2BxgKDm+DI6lw2XMxk42oBMWSZGflA9FDFtQwaPT7bZh30
8qMQtteMYJPumFFTSuMlgX2CTtkFS67JSBZt7Ixesot/vep/1noZ/h5XWn+gV0IhI/uDSd714eVU
zOCJH9U7C6VevG7VGlW8RKORnPu8fBNm1qEijgUnJmZQlQ+1GyvLDSWNBnI8Yhh0f9x6qd/qrQ7H
0qHm/WVTbTWHgUNwXCsW5Kw4KKasruKeUPpKBJQBcy+IgO5W1lewUbveAm0gYYqx7IfZBNfRgrgg
ipFNkYgVtTSD9S4CQUP29DmW7/VthVw5ey+PYdwW0h09ckRfIqDp5A+DH8QelZ/QnmurKyScMMB2
232ZYB/gGMYYLHl4zlnzs/KTwXaiFMKWfiMeC8RQOJAQYnWpV2+9kIX7fPGkh3j/fBqvGVxhhWVf
ZbuJriZaMXMhAWuobhKmAYbG9vHHhBtkAtKnmAtMG/L56m794kd+lK38rJx3ipv2j5YNkJzJ3mr7
2XcFM4odByre+wi6qB8efzi9MmwJ2KGmDjZ1lncmikZzH+GSHZuQJwaqGFIs4s6A7iqNg24TQS7r
3Pw43TgWmNNwY2xyoUQqHf61olqKg9MVhEgovzP4+bfrRdYXXLqGZAg/F5xbiO1PSer//MlDxlo6
9EfvDFwruWC2qS9+2rBscu9UkrCZeMbPn7jFVcygN8A9g5Kup654o33hRuz4il9w6J3cr+1sVzOg
XJWBgequnnM+fV2o5QfXMXi2wTPMdHYl/glJ/1o9aGRZXIU/62CiwRwdI3em3E9zd2TyNwN+a2Im
QPIcPE+1XwWZi3Uj8tjvBbQaFc31IclXGImhYwhBR5kiSzr/RFqJ6O4GtQLJ2WiMdMUw60bs7z75
U9dT+W/2JLkNJrYmhHP+y+Tv6gfjpcHvNJizlpB31EEQwpJR/3+WoTsJiWrHmy4xGHmG4wwhz0zs
4wjniEUNsB2rlwQjvleO6owO0QYd9frbtctIqWoDfR6XPEIKUQ6H9ZTftDzM7XPZAW9ItSwDXvvG
4pUSmGlvgnOV+yVG6DfJBzCFkHGdkQY2oeTbh9GfhZ9AW3yIkEXyzfKtCDM4WGldPzkyDWY4sqCm
SRCOTgx7OWAVstXdglZehwBWQ6Sds/S7j0FZefh4/yndByIGQBSOBfPaPQMnTcXT9KUTcKvHTTEX
Eu1qnrMGgE9vERPFvdMfU7Y9uqXGb1PC4bsYw8isvfR6MZ+WcbNZdUdXTnV8SzCc5BP+HV6OViL7
JBCwME5UiDIIGNFiMon6e3BXzfj8fP1pF2o2nzHNuFu4KPBTOgkbOYwhEDaHpy3mxCG6sHH5vVz4
YZ73q9zXZ2JiW1ExRN92PHMgofuJSl4Hu4pmhUF1a9RbLCk9rXrIYArDG3cDIQlac8tBbXT4mjXR
A3JdQrf5/zNWDp0G/LTGqillxoNSscik0RJNnFW9WWVcLWqxAz+54YpWpIiD4LzvbAzRwNGNQLNB
t+kMTE7O1MZANEUI2zmcCWEIU7j7ovW3tDf2RP7HW5boCWV6CiRpyosMzYD9dqcKOKGfj/sqkxt+
b82CFVObv2w2OtG0FjJTCMpsZ6HheeTawgFUiMsqvqafDHHjKhG8ASWGPyENNy9R3i+y02BCVInw
GNAnn8Pv+h8NUeqyqZdBNcmazw9iPMLEp8Ma3WvKqkJGaD1zgPNkkfEHzQM9JcS3ZsUYcwCre8He
oV/kx9kD8zv7O/p+lIctN5IpmQSEBlZdoHE3qHn6Ublii71gMSvZKjfF3LPERTcBRv6UfUeqWeVX
229RBmRGm6PT8rt7MXxhhwCir0r6na3dv2f6TH55ss2puS4xekIXVwOW4FAZkGP0wU0WB2YOyKCD
SAVn7dmAAMtYuxjboqL7drk4zBVgDiMqlEW66oblr2kB9LEpzIpe3q7y3JBDNkI5eDnsU7OjXmaz
8RiTdyjG+tK5gkHgwPuOx8mARf+8vd7m0ZAGKQbrXmFk8NHrQn2ezN9a4b11CfuF3yriZUD0uQ1L
yWpkzQT9Ns7CJzhoGEgRQGiMzlX3XTVBT4ZjZ588rLdPCXnn36ZdOw+L1woxwb88MKyOQ81pgFZq
hTXm6diV7sT8pLPycqCoAcBUrpgy5iM86jBcl82KPEmIQnO9EezXB4lkzt6j4l5jjCdX5IpuCsxv
YFddK34IunrgkxttNRPEyC4kwhIa4F41FMbmnGZKqWBdN8hFoFfNQPtsbOy/SVyiizXBhBo4eKYE
w4lRPjMfPDDRB3J+NcpY8bBW/Nwxz7EicKspzBwRQxADI3nLWihDrH4UpXuteHLzEbN8bAkAncQo
tAsSLMR1WesmFDRCZvNum80jMjL1cwnBI1ceicLlmhRu485VHbCuFr76d6PYyxEAuV+FZl8Xhe8h
AwH4HkWFRkOa3jvqUB3vqUY7XeVlQOtre7qlAeYgR+fDkzBO5LAn00TlaLLvgerXLSVawGxg4r2N
6KJWsunna20ThYRzLx+i1k1fkshaY9QqbzrohIYqMGZQE+XsE6qqPXsvd4gvLjxnfWVNLQH4UEIV
pZNVfWTIPCuehYspvcOK0f0CEIPZleld1CB0TwCxCN+S9yN1WIu+i4YpDf9V8kbVDylUnCQjKAWv
T+2go4TgsZpzcrU1XA/rA0EfFWxiJvAf7QssOMv5QVo4SztdVxeOm75FNlUMj81csI30WitQ3hYh
oqAGWq3MFPhSLMWRWmaNzuw3g1Ve1s7fg7o+/kP+McJwxVekkw8gk1dSVt/VoA0Dgb6hP2DJBwsd
NBSNMI+D4k4pqW2+CnH79d71mR4T/VRyi0XMGjahoI0ttUJfElLP/D3lk+7+PZ0eTyZ6pv2jfNKE
TaAql+mZ91yGnWm9md/aaTw6aTY7ywOjeOgUTwmkZiNX90BiMBc+dMHY6ZzLrHEK8t5Enk/JWu09
ZRoHRGAEHeNIO0t1GtuM0dHZkZpO5nyHoKKmn9CIHeGaQ1dN3CZGEdaN82FMfVNOw3xfg45Lpx43
zlTobi8tIs7DCmaWiwP7nZlVe3oyh9lfyR51Dg/6jac2rNPaSgHEsmSmjmRcmvUPecOatxcUPvid
S7jrZa9Lt1+XGS86FD6qHdFO2BfGFtuEe5jlCr6MwFkEhcINP9PWMpOiZWZdb8q00RkuQwMaNOse
f71syW+viqJbZGVecKTyuH2LLrNXDce0OMfOe7fYWgc8RMc6325Jmq27lo2LlApzdNSEGqo4A/1f
k0tDUchitnfGFngNOzNUwhIX5emiCnRU3DwZnVUR5hAFpnafRZZTUNSsO1EcKT2fLCtuBhzb39ZN
RNwWRKcZ/wj4vhGyBqwq+vUlYhs4Dys0HxO+LEKAy/l2Iiws+s9NNhbaneW8w+YV5VVpl3NvhSgS
FY94ugSt9/+ZFxD2f0pty+GaFZ4y4187G8qZWc0LaMxrt+QzjGKKSjCkUS5zvtjaCUHojsjYwale
IdS+SBcr9cRqOpx+vNKsFBr4Wm6NpJcRJuxOo1SeyZPOKACT3q1ngwEcg1TlEpYPgLEiuMlykBRE
/kx8e1HWRdLlPdjUPhSZ6nJBntL0Fmz0Y2Pi8Ff/FvQ4BdBEe+b2yiM8ALla4T3BfoweitA4/+vX
7OzOuU2ePYplQI4dA4e8Xmo3OVOblp4lvN83fFNgofX69607jMIwtr/ufyrLyAce77L25U7e/Vkz
MkmX3L4rifg1KjCcn5N2+V3VJV28GD3gzyCguTBa5ArGH6AonxjOPFiHIg3+8Ly6hn/DISTgQ0Vv
5o87gfLi/au7tZ+/rUEF1OVlsa3xSqYs3t5TPYJgonaL450BkTWg6kHlD/fyw0TjCbRSiL6jYYe1
GxCduaqEtIIouS+E4xGPUW3tuJ0wZHWMsWS8FZLECUI2yCEw3WqGkAVDfcLh365XjmIxbbmUNTZB
XaoY6CF9aP8Q1c+sC6oEQY02Oi5YR0CeUk/BusLwtw6Z7yqMDyGBPC4THoI+UeFrMVBmvZ2itFDL
ZbFzE7gjiZ6lYgbi/O4Brr33ETzLmjV/VYikI4tkRgZWLJjdSGOZvH/f6VZ3v3v+EOD7wpPibjmm
LPp9K+RXNqC2JZrVdpyykw5i9IW/ytIyv4Omc2cmLzrlsVDbafbcnY5s5XGbmSOfx0YxWkIKnuNm
wX0CjZOTDOHsuO1O/FR3v0yrPsCNoxKslSRkr6RCjmll4zlOp9+IR8ygGMf9X69L+gjZ7mreZxmb
zd7rOO/yo63lHucCIULLiXI0adrgbVigne+lyte1MEI+PZLWlQnxwfnitqchMFazC/v2kS/HQaXI
Nc1H5VYqYgM67I+PwM3laICMlZSr8YKIwDzdvexTOSyKiNmtJJTrO7L9ZOBUHzzjYuzZn/rIVnhv
08jrPeM1wdSPQgNsubpOaqXeUXN0vcd2C3oCqGKm0NxqGdlZbSBZqKB5PjSdEGUQL2lfJ89orUdb
ryzaAQKK/DeeyKqPqRE0abocvUhBJOG9MwZGMrgA0nsRm2DvdXgdpfBFxOUxOi4p+N+OmIbRAAZO
dT/h2wyLcbIYqer5FYD3Ti3ZeVtIJpUJ4ApsSuosu24IEsAmKGdorIqnXaums58rVps+Yn1nzkNm
dpd0AQgb1KAtxTCJUXMM9w2MIP5Sv+G6hofhT56dsA5xWRJUganYbtdgN8mZQWn7tGNGJAMgznjp
CR3nqHxNySgzlbfREHNq+fqXE8n/BGIV0Bxe7I0YZ4bnRuumhaZ0E0YRikpPX0TGI/N1KvqTkc66
+BQ3dn+zds/7e1UnCn86yVBt3sPeDOS6u66RxFoHfuxfbysp4Ty/RuDNi4Fme0WlO/QGNvwuz3aD
nvoc8N7l2aDZHpbijysFk1pjp0+ca9OlC6EFGoQRQgXSuruXnMbZxT+8cH4/PV07CIM0gDPog/gu
XDSiWXQ4MRUCS6IyES38BheHGoWELgpUk08mFr3h+x0ySDEO+X65INEp+hhj4xMLLV8XOOX+Ezz0
BFAXmfTB6Iko0svFosyQDSvfFA7k+/sDSHwzQtaoPQjct4KEmoKcx6Rd6k16SzVTwX0z9ofGlNR6
xGib10jEcccOfOSBnaA9ErCylbTw3r78sxtg+XXo564JsYBUFQLcQMaI8YivqF+MjkNOvcs29U2n
nT3+UvE/TR+FsG1KzJ0aCMMblKFPIEPJBXKNFiuXTmXuW4BZomxA/k18yBEqYrgR5dBVv+VSBOxb
qohDHYompx4ILHCjp1xmKJk4cNBdCkU5arjx1Aedp955DKlukNk0QnkB2yBvec3sLHr/HbXCzDDu
+J1JJ41ps6xutb3TlX4L0VHwlQ3h5pHfBKRVHy9o4laHYW4I/5dqIAmq0PiNTPDI716rjOLa4MmY
JPuOe1SLj/x9RuC2Dc3+FHe/NZT5Z/X3bnxkajU3B4TFfwHLqhUxd6Dqu/c0EZ/FOAHEzNXbEXX/
e/3K/x/DKu0XeOhxa4CFjtzMhuL5KVTgZ/VF63y43pmcbmtzow7pcBxEGJkY28TF10xokNzF4WY4
x43YdB4Fumiq67zMgMzSRTXBgLM/D00O2xZOdmFhrVL0CRFSQXKyuJ4+RdEkmwBI1wWOu/aqURch
ak+HYX7IiJjKqRFSE/HkQzhboa5C9gdRmdaZMAxp5eAfUd6pP8prwFNGOGOfXCw88FSvt4aIkzcN
bU0qHtiLq9UlPK/J487X9WKo9hujWJUjt7qqgOOgJxQLjVwkk3Dx69oIw4O0K4pEGGsgLVRdSVtz
7ACBbGkaQ9VUL4zEYoFfuKsbMtbPlVTrp964gSIU/0v2jU/NQjxCSTH8Wfng8P5a0tzlFwcgp0En
KvIWWbSNJCzn2uY7IQtVS5ePU8m82WmWisUU1O8Qce+4OwoTrdpVfkMV9a6noqmQdnRgvrB+HaOX
6T2+vBcftlYRwOv1ZlhLIsnhYDNjgH+KTLN95ZDtrXBBVmVMQ5mIOkSpzw3rnqzMfEaGDtfZzG+T
9EYhyBhtEPZGyFtFsQ80BLikDJjJntVF0Vk+UMR6IIkAJihQYRIqcY3n2+sYLDAqEGIks/M5njTr
H0QZIe7pkNIsD+BAzv4RbgDmxKAbCI7v/sXOXwETi/LoxYgVQrU5lf5R5n+odGhmTwEj+r/Wl3EQ
tUCHod6vn9gy3g9FtE+NTq/z1QwzbkSaav/Q5m3hsuNvmGJjb0/Svbzyt/8az+KijHau1QciBOrl
g8K4XY//f4Zw0V3eHKUmHxUq4uYT4f4RWv5+NYeNjGZo6cmL0XWli6QBefdRJHvzm29Wef0WVfPV
FgvDYdkM/pYWcrZZru8Pe9TCdtiU7ubefkl1+AbGIjq+xt1k4XGhIYy8t7Xxdkd3jiaMAXMiTLlw
4td9feq5kEFXG98UGfxRGmKn6MY1+aUCJJ2MZO4zzeSrS5CvOS8fnUAV/yJ+Te0EpCI68jifu99B
pmot2xVZ/SrbvgaO3DnP8yaKKzXLp+IhS9HasEGr9w65dupzmqo3IKHlco8fwWcI2tFBJV7I4bgf
bDamHWq2qojK2tYxcdZxlhCwN3uONre5d+0fY8B/S93vN1jT99d2e/CznBh4wiOoB3YhYvWsB51D
WZPepQ6bzirALStyMRPKYOx3J/DSlnecb8MAakKHndNqluI2d+MzJu9URwYLRbGK6YbgB+xfav47
nu8RUgQdBWYNgCmR5bzx6oH/68PghJ+K+7OOdx1ULEurqSnN6YbzzR1u4FLNv4/QJPYi8Pk9c5F+
3qZ4VRLl04IRwkxsJOcGdct9dA3ec3V1Gu53bV+2p1Qzv6PXhjPj80kbnvr8dsti03fa4bvv/A4k
rrrJOmHJvw/CLmXzJyFyOEUaZiFsIts5aXTrAGXz0o547czSXsMI1l+MeFLONa8XsYe/yDplhfo5
GXSpjt4ZFBjkoRBqC0vh8t1nsKaZDzRM+5XHLcE7xGVTk2y9odB0NJ6YZQzU+6uSgFzN9Yfverae
5d8fDNsWYweHsbBENYdmQQSfwjJR1f0Bf9X1rP7cLQhmlTxChObSJ2QG5XvPiLWptQYipbXIG182
TEw/QzUnmJR/YE6DdbcnrmHRolcHiIyVTXXeHjhKfSmgxilYPOIqsuVC8wHatoA2RkDeJ4hyZZRW
0jF+YUkVTb5epwpDbWmo+YIlfXx4cUXxRRE2R0Hn0DypAdvVz4k3P6nh2Q0eEfHstgxetAe5SATx
cC8OeHBrKw7ISOT1Yt6EZddhARnlTuVFZGCx2IFKep5jGrq+a1K855zbw4E6ovEOnKYrQ+HT9yvk
e1PDYCBw7ot1qRWyJVw/Hu2z+HXp3K5f8/EAmToEofVzZKs4VvPK7B3atrulv+80hbRDHOd5PUjZ
TyP17qbqIi3BTRHOUebC4yWVzUvehzXaFs+7HFx37HPQBeHwlUQLH/bQfzAGEBn28/r+rV7cXC35
XEf5hc2kCmUyroCIUIF4nysO5eFaHkeqzn+MtwWV/L1HsoXuu7TGdGerWdSpesZnuMbqozJiKq1N
lNUbKQsJdtRvYfQgUqGoklKvgoTHLt6W2APXWjcWrSPj4vzpm4RNkl2nQi785rNwJb3v4QBa5Uk4
wdb03OM2EVdL3PmevllnvfbcO08GQoYOSLAiTb+ICEFnDtOHNUPRHxrkZtW2H4Jqj2qojMAnVZ7w
T07NUd9Kg/UWwj2bJLxnODodd+UATh4I/gX/fXbIIYRnq5Uh7aTwgUZsdHlDC83erZUEBACz7uWa
iB4/mo94nKmbGUQHAc257y9MECqPDpRypS+oYJCMO5pK7OX70nMBhEvyXO81iOpaaOhw2JHsF/yL
Tp6w1A9Kzh3pFDDMsYA1Pc8VstT/6D2QpGGZ5LZxnJUVOGB+oJRw0/X71mUH7KKjtOcKvBw55aSZ
wy7ZFPxwagRb9amDNEIrVWyd8k7JfXZ0CDV+kJK2v21c3SE1VttD9vy8tU+xLzzy6S4nwdV4vOa7
JU+Lm1pKq+th509apPorYkdAUsoYb/TAlGtjB3vbJ+ZEcRIQNepISnQEPyLA2fZ3QLu4xJmAua/0
UOK8DwHaF1r5SddiBFKAJg/KDnXfKOBdt68cmXuuxgVlIBH1ws+uhP2mdGAK3ZA5pXn52GKkGOUW
+WdAwIBBhTza88S0hhDnidfMlWrYqyZdCa2Myux4+2YrtbGI/UvDiWNYw5VCDo7OldEkQTAzV2R0
OTZnRnGQiodB80ylIn4f+1y49e4zqhj8auJj+we7Z7MTVs8VHfFIhXiv8rzBgI12OcfF3AVM3EFi
Oiw0SbzzMvi3T1N4FLtympIXedQ1JkTG3EJ6R2Ds376ZhjA/B1q/fZK3hzfsjy8k219eThCIodM+
bHZnVk+6Bcdvay/UtiYESx9FU6Sj47JK+F2A3PuZ6gkL0p72SrhNakA4fb/c97/PPfm4w1gGO5cD
MqSlcUeqm9hwRTKjbI/AJBAxCUa3YEfLrA90UKVzr3JLhjCvvPbdBYMTyU8moIkqyJI6ILYxFR5J
2aWD32sECNuFi7TGY/XVfTkS7omQbaKZ5CS8u1nERlDAe/Z/b7V9GNEPCbzyTzggN6whqh++maSp
XAsib7g1HVYJSeKL2K3yT2oinZ7RYxrghCHJBt1XYzkSBAuQFo3Ugv3FX6htlp3CgCXkxCDwhfrQ
h3S8yr4GnFoDD2wl9412IPEb4nf5jR2g2fWmIU52r2QZK8zwgVg21XzoHWUxlTMQcje1cDm+Hqpz
bc0etR/wf3gOSf9jiePJoh4PTXvnHlJgpIsiup/G2mKfX5VQdjvNiDQx6WKx0NsI5XH+Cs8m9eO/
czJc7nOWxr8slxAgzYNPBR5TXJeRz9M95MueikvSASS8zJKtAq+2wTTQOAPslTeZgxWrfJ8PTYqX
6uK/abJ+Sep4CkGHaWmBN+q5sZShiZcqgizE5obBzf1w1dLlI8Cz0badrQmpEhJYMavEhqWZr2mD
yhQa5fpa9BB3ToNgLvkjFEaWnB/ii3fNgmdjhlKgiX3ke35zc21NQW3/XdJJC9xOs169e8Nrea3F
cEcJqPvsXgLUhrgz8peoOOrBJBYKB/0GoUs84Xo0AIYxLPxRaDhIGJFAdM5TsUGssXzUE9bGuGfo
rnEKzr81CRP586AkuwckBlDHlpiunZ+075TlSXWq8oDC3FgJI2hoYTdS2letBvYy4pwXx58nyqxA
UDBuCyRNLR6EJAfs6XTlpJEaEvE2R8WVNxsi/Hdx5MqL04erNMyEDzvJVWvuGV6KEcVinxMAsB+4
Ql5qA51XDwk4UiUBrakE/+2P3Vtc8mjMd5bZ5OY1rQKKRDSFUuRZ9OrC2pNV/+G2E5DVS/AcktxB
AO7QbRT15pE7LrAdpI1Ux5/M58XSykFDRGkRATsTWa9dZRjDVJ14IPewFG/G
`protect end_protected
