`include "sample_tests1.vh"
